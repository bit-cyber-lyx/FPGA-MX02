// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.11.0.396.4
// Netlist written on Thu Feb 25 11:55:51 2021
//
// Verilog Description of module system_top
//

module system_top (clk, rst_n, key, led, rgb_led1, rgb_led2, en, 
            one_wire, rs232_rx, rs232_tx, piano_out, oled_csn, oled_rst, 
            oled_dcn, oled_clk, oled_dat) /* synthesis syn_module_defined=1 */ ;   // g:/fpga/mxo2/system/project/system_top.v(1[8:18])
    input clk;   // g:/fpga/mxo2/system/project/system_top.v(2[15:18])
    input rst_n;   // g:/fpga/mxo2/system/project/system_top.v(3[15:20])
    input [2:0]key;   // g:/fpga/mxo2/system/project/system_top.v(5[29:32])
    output [6:0]led;   // g:/fpga/mxo2/system/project/system_top.v(6[29:32])
    output [2:0]rgb_led1;   // g:/fpga/mxo2/system/project/system_top.v(7[29:37])
    output [2:0]rgb_led2;   // g:/fpga/mxo2/system/project/system_top.v(8[29:37])
    output en;   // g:/fpga/mxo2/system/project/system_top.v(9[29:31])
    inout one_wire;   // g:/fpga/mxo2/system/project/system_top.v(11[18:26])
    input rs232_rx;   // g:/fpga/mxo2/system/project/system_top.v(13[29:37])
    output rs232_tx;   // g:/fpga/mxo2/system/project/system_top.v(14[29:37])
    output piano_out;   // g:/fpga/mxo2/system/project/system_top.v(16[29:38])
    output oled_csn;   // g:/fpga/mxo2/system/project/system_top.v(18[18:26])
    output oled_rst;   // g:/fpga/mxo2/system/project/system_top.v(19[17:25])
    output oled_dcn;   // g:/fpga/mxo2/system/project/system_top.v(20[17:25])
    output oled_clk;   // g:/fpga/mxo2/system/project/system_top.v(21[17:25])
    output oled_dat;   // g:/fpga/mxo2/system/project/system_top.v(22[17:25])
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // g:/fpga/mxo2/system/project/system_top.v(2[15:18])
    wire clk_1mhz /* synthesis is_clock=1, SET_AS_NETWORK=\DS18B20Z_inst/clk_1mhz */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(18[9:17])
    
    wire GND_net, VCC_net, rst_n_c, key_c_2, key_c_1, key_c_0, rgb_led2_c, 
        en_c, rs232_rx_c, rs232_tx_c, piano_out_c, oled_csn_c, oled_rst_c, 
        oled_dcn_c, oled_clk_c, oled_dat_c;
    wire [11:0]tamp_data;   // g:/fpga/mxo2/system/project/system_top.v(25[21:30])
    wire [23:0]time_data;   // g:/fpga/mxo2/system/project/system_top.v(26[21:30])
    
    wire flag;
    wire [9:0]data_length;   // g:/fpga/mxo2/system/project/system_top.v(83[14:25])
    wire [959:0]data_buffer;   // g:/fpga/mxo2/system/project/system_top.v(84[14:25])
    wire [2:0]cnt_init;   // g:/fpga/mxo2/system/project/ds18b20z.v(37[13:21])
    wire [2:0]cnt_read;   // g:/fpga/mxo2/system/project/ds18b20z.v(41[13:21])
    wire [2:0]state;   // g:/fpga/mxo2/system/project/ds18b20z.v(44[14:19])
    wire [8:0]data_out;   // g:/fpga/mxo2/system/project/ds18b20z.v(46[20:28])
    wire [19:0]num_delay_19__N_369;
    wire [2:0]state_back_2__N_261;
    
    wire one_wire_N_501;
    wire [3:0]tamp_out_11__N_478;
    
    wire tamp_out_11__N_483, tamp_out_11__N_489, tamp_out_11__N_495;
    wire [15:0]cnt_adj_5212;   // g:/fpga/mxo2/system/project/oled12832.v(28[36:39])
    
    wire n438, n439, n578, n579, n580, n581, n582, n583, n584, 
        n585, n718, n719, n720, n721, n722, n723, n724, n725, 
        n863, n864, n865, n998, n999, n1138, n1139, n1140, n1141, 
        n1142, n1143, n1144, n1145, n1278, n1279, n1280, n1281, 
        n1282, n1283, n1284, n1285, n1354, n1355, n1356, n1357, 
        n1358, n1359, n1423, n1424, n1425, ready, n26793, n29, 
        n25772, one_wire_out, n15, n16602, n5709;
    wire [9:0]data_length_reg;   // g:/fpga/mxo2/system/project/beeper_control.v(22[21:36])
    
    wire n15_adj_5200, n12, n22685, n23656, clk_c_enable_684, n5151, 
        n4, n20945, n23969, n23972, n23966, n23974, n23973, n23971, 
        n23970, n23967, clk_c_enable_688, n25484, n25453, clk_c_enable_659, 
        clk_c_enable_1399, n15_adj_5201, clk_c_enable_1439, clk_c_enable_931, 
        n37, n28, n25806, n25618, n25765, clk_c_enable_1437, n25751, 
        clk_c_enable_132, n25742, n25607, clk_c_enable_686, clk_c_enable_1433, 
        n50, n25824, n25774, n25773, n26780, n25706, n16451, n25857, 
        clk_c_enable_117, n25689, n25826, n25685, n25825, n25808, 
        n25807;
    
    VHI i22683 (.Z(VCC_net));
    LUT4 mux_123_Mux_0_i31_then_4_lut (.A(cnt_adj_5212[4]), .B(cnt_adj_5212[3]), 
         .C(cnt_adj_5212[2]), .D(cnt_adj_5212[0]), .Z(n25825)) /* synthesis lut_function=(!(A (C+(D))+!A (B (C (D))+!B (C)))) */ ;
    defparam mux_123_Mux_0_i31_then_4_lut.init = 16'h054f;
    LUT4 mux_123_Mux_0_i31_else_4_lut (.A(cnt_adj_5212[4]), .B(cnt_adj_5212[3]), 
         .C(cnt_adj_5212[2]), .D(cnt_adj_5212[0]), .Z(n25824)) /* synthesis lut_function=(!(A (B (D)+!B !(C+!(D)))+!A (B (C)+!B !(C (D))))) */ ;
    defparam mux_123_Mux_0_i31_else_4_lut.init = 16'h34ae;
    ROM128X1A mux_415_Mux_55 (.AD0(n25685), .AD1(n1359), .AD2(n1358), 
            .AD3(n1357), .AD4(n1356), .AD5(n1355), .AD6(n1354), .DO0(n439)) /* synthesis initstate=0x0000000000003C3CFE307C20383C1038 */ ;
    defparam mux_415_Mux_55.initval = 128'h0000000000003C3CFE307C20383C1038;
    ROM128X1A mux_415_Mux_47 (.AD0(n25685), .AD1(n1359), .AD2(n1358), 
            .AD3(n1357), .AD4(n1356), .AD5(n1355), .AD6(n1354), .DO0(n578)) /* synthesis initstate=0x000000000000623C307C662438601042 */ ;
    defparam mux_415_Mux_47.initval = 128'h000000000000623C307C662438601042;
    ROM128X1A mux_415_Mux_28 (.AD0(n25685), .AD1(n1359), .AD2(n1358), 
            .AD3(n1357), .AD4(n1356), .AD5(n1355), .AD6(n1354), .DO0(n863)) /* synthesis initstate=0x000000003800083C0C3C3C203C7E1038 */ ;
    defparam mux_415_Mux_28.initval = 128'h000000003800083C0C3C3C203C7E1038;
    ROM128X1A mux_415_Mux_19 (.AD0(n25685), .AD1(n1359), .AD2(n1358), 
            .AD3(n1357), .AD4(n1356), .AD5(n1355), .AD6(n1354), .DO0(n1138)) /* synthesis initstate=0x000000000000231C103E332418201843 */ ;
    defparam mux_415_Mux_19.initval = 128'h000000000000231C103E332418201843;
    ROM128X1A mux_415_Mux_0 (.AD0(n25685), .AD1(n1359), .AD2(n1358), .AD3(n1357), 
            .AD4(n1356), .AD5(n1355), .AD6(n1354), .DO0(n1425)) /* synthesis initstate=0x000000003C0008630C66332026061826 */ ;
    defparam mux_415_Mux_0.initval = 128'h000000003C0008630C66332026061826;
    PFUMX i30 (.BLUT(n15_adj_5200), .ALUT(n12), .C0(cnt_adj_5212[3]), 
          .Z(n22685));
    ROM128X1A mux_415_Mux_7 (.AD0(n25685), .AD1(n1359), .AD2(n1358), .AD3(n1357), 
            .AD4(n1356), .AD5(n1355), .AD6(n1354), .DO0(n1282)) /* synthesis initstate=0x00000000DB0010630843402360181843 */ ;
    defparam mux_415_Mux_7.initval = 128'h00000000DB0010630843402360181843;
    ROM128X1A mux_415_Mux_2 (.AD0(n25685), .AD1(n1359), .AD2(n1358), .AD3(n1357), 
            .AD4(n1356), .AD5(n1355), .AD6(n1354), .DO0(n1423)) /* synthesis initstate=0x000000001C00043E043C1E201C7E181C */ ;
    defparam mux_415_Mux_2.initval = 128'h000000001C00043E043C1E201C7E181C;
    VLO i1 (.Z(GND_net));
    PFUMX i21094 (.BLUT(n23969), .ALUT(n23970), .C0(cnt_adj_5212[4]), 
          .Z(n23971));
    PFUMX i21097 (.BLUT(n23972), .ALUT(n23973), .C0(cnt_adj_5212[4]), 
          .Z(n23974));
    ROM128X1A mux_415_Mux_54 (.AD0(n25685), .AD1(n1359), .AD2(n1358), 
            .AD3(n1357), .AD4(n1356), .AD5(n1355), .AD6(n1354), .DO0(n438)) /* synthesis initstate=0x0000000004003C3CFE307C207C7C103C */ ;
    defparam mux_415_Mux_54.initval = 128'h0000000004003C3CFE307C207C7C103C;
    IB rs232_rx_pad (.I(rs232_rx), .O(rs232_rx_c));   // g:/fpga/mxo2/system/project/system_top.v(13[29:37])
    IB key_pad_0 (.I(key[0]), .O(key_c_0));   // g:/fpga/mxo2/system/project/system_top.v(5[29:32])
    IB key_pad_1 (.I(key[1]), .O(key_c_1));   // g:/fpga/mxo2/system/project/system_top.v(5[29:32])
    IB key_pad_2 (.I(key[2]), .O(key_c_2));   // g:/fpga/mxo2/system/project/system_top.v(5[29:32])
    IB rst_n_pad (.I(rst_n), .O(rst_n_c));   // g:/fpga/mxo2/system/project/system_top.v(3[15:20])
    IB clk_pad (.I(clk), .O(clk_c));   // g:/fpga/mxo2/system/project/system_top.v(2[15:18])
    OB oled_dat_pad (.I(oled_dat_c), .O(oled_dat));   // g:/fpga/mxo2/system/project/system_top.v(22[17:25])
    OB oled_clk_pad (.I(oled_clk_c), .O(oled_clk));   // g:/fpga/mxo2/system/project/system_top.v(21[17:25])
    OB oled_dcn_pad (.I(oled_dcn_c), .O(oled_dcn));   // g:/fpga/mxo2/system/project/system_top.v(20[17:25])
    OB oled_rst_pad (.I(oled_rst_c), .O(oled_rst));   // g:/fpga/mxo2/system/project/system_top.v(19[17:25])
    OB oled_csn_pad (.I(oled_csn_c), .O(oled_csn));   // g:/fpga/mxo2/system/project/system_top.v(18[18:26])
    OB piano_out_pad (.I(piano_out_c), .O(piano_out));   // g:/fpga/mxo2/system/project/system_top.v(16[29:38])
    OB rs232_tx_pad (.I(rs232_tx_c), .O(rs232_tx));   // g:/fpga/mxo2/system/project/system_top.v(14[29:37])
    OB en_pad (.I(en_c), .O(en));   // g:/fpga/mxo2/system/project/system_top.v(9[29:31])
    OB rgb_led2_pad_0 (.I(rgb_led2_c), .O(rgb_led2[0]));   // g:/fpga/mxo2/system/project/system_top.v(8[29:37])
    TSALL TSALL_INST (.TSALL(GND_net));
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    ROM128X1A mux_415_Mux_46 (.AD0(n25685), .AD1(n1359), .AD2(n1358), 
            .AD3(n1357), .AD4(n1356), .AD5(n1355), .AD6(n1354), .DO0(n579)) /* synthesis initstate=0x0000000030004266203C3E2C60601042 */ ;
    defparam mux_415_Mux_46.initval = 128'h0000000030004266203C3E2C60601042;
    ROM128X1A mux_415_Mux_45 (.AD0(n25685), .AD1(n1359), .AD2(n1358), 
            .AD3(n1357), .AD4(n1356), .AD5(n1355), .AD6(n1354), .DO0(n580)) /* synthesis initstate=0x0000000068004266200C1A2840401042 */ ;
    defparam mux_415_Mux_45.initval = 128'h0000000068004266200C1A2840401042;
    ROM128X1A mux_415_Mux_44 (.AD0(n25685), .AD1(n1359), .AD2(n1358), 
            .AD3(n1357), .AD4(n1356), .AD5(n1355), .AD6(n1354), .DO0(n581)) /* synthesis initstate=0x0000000040004242200C023840401042 */ ;
    defparam mux_415_Mux_44.initval = 128'h0000000040004242200C023840401042;
    ROM128X1A mux_415_Mux_43 (.AD0(n25685), .AD1(n1359), .AD2(n1358), 
            .AD3(n1357), .AD4(n1356), .AD5(n1355), .AD6(n1354), .DO0(n582)) /* synthesis initstate=0x00000000041842426008063040401442 */ ;
    defparam mux_415_Mux_43.initval = 128'h00000000041842426008063040401442;
    ROM128X1A mux_415_Mux_42 (.AD0(n25685), .AD1(n1359), .AD2(n1358), 
            .AD3(n1357), .AD4(n1356), .AD5(n1355), .AD6(n1354), .DO0(n583)) /* synthesis initstate=0x00000000041842424018043042421446 */ ;
    defparam mux_415_Mux_42.initval = 128'h00000000041842424018043042421446;
    ROM128X1A mux_415_Mux_41 (.AD0(n25685), .AD1(n1359), .AD2(n1358), 
            .AD3(n1357), .AD4(n1356), .AD5(n1355), .AD6(n1354), .DO0(n584)) /* synthesis initstate=0x00000000041862424018043046461866 */ ;
    defparam mux_415_Mux_41.initval = 128'h00000000041862424018043046461866;
    ROM128X1A mux_415_Mux_40 (.AD0(n25685), .AD1(n1359), .AD2(n1358), 
            .AD3(n1357), .AD4(n1356), .AD5(n1355), .AD6(n1354), .DO0(n585)) /* synthesis initstate=0x0000000004186666C010042064661864 */ ;
    defparam mux_415_Mux_40.initval = 128'h0000000004186666C010042064661864;
    ROM128X1A mux_415_Mux_39 (.AD0(n25685), .AD1(n1359), .AD2(n1358), 
            .AD3(n1357), .AD4(n1356), .AD5(n1355), .AD6(n1354), .DO0(n718)) /* synthesis initstate=0x000000007418184208C6422046041046 */ ;
    defparam mux_415_Mux_39.initval = 128'h000000007418184208C6422046041046;
    ROM128X1A mux_415_Mux_38 (.AD0(n25685), .AD1(n1359), .AD2(n1358), 
            .AD3(n1357), .AD4(n1356), .AD5(n1355), .AD6(n1354), .DO0(n719)) /* synthesis initstate=0x000000005418104208C242FF420C1046 */ ;
    defparam mux_415_Mux_38.initval = 128'h000000005418104208C242FF420C1046;
    ROM128X1A mux_415_Mux_37 (.AD0(n25685), .AD1(n1359), .AD2(n1358), 
            .AD3(n1357), .AD4(n1356), .AD5(n1355), .AD6(n1354), .DO0(n720)) /* synthesis initstate=0x00000000D218104218C242FF40081042 */ ;
    defparam mux_415_Mux_37.initval = 128'h00000000D218104218C242FF40081042;
    ROM128X1A mux_415_Mux_36 (.AD0(n25685), .AD1(n1359), .AD2(n1358), 
            .AD3(n1357), .AD4(n1356), .AD5(n1355), .AD6(n1354), .DO0(n721)) /* synthesis initstate=0x00000000DB18304218C240FF40181042 */ ;
    defparam mux_415_Mux_36.initval = 128'h00000000DB18304218C240FF40181042;
    ROM128X1A mux_415_Mux_35 (.AD0(n25685), .AD1(n1359), .AD2(n1358), 
            .AD3(n1357), .AD4(n1356), .AD5(n1355), .AD6(n1354), .DO0(n722)) /* synthesis initstate=0x00000000DB00304210C2402240101042 */ ;
    defparam mux_415_Mux_35.initval = 128'h00000000DB00304210C2402240101042;
    ROM128X1A mux_415_Mux_34 (.AD0(n25685), .AD1(n1359), .AD2(n1358), 
            .AD3(n1357), .AD4(n1356), .AD5(n1355), .AD6(n1354), .DO0(n723)) /* synthesis initstate=0x000000009A003C4610C2402240101042 */ ;
    defparam mux_415_Mux_34.initval = 128'h000000009A003C4610C2402240101042;
    ROM128X1A mux_415_Mux_33 (.AD0(n25685), .AD1(n1359), .AD2(n1358), 
            .AD3(n1357), .AD4(n1356), .AD5(n1355), .AD6(n1354), .DO0(n724)) /* synthesis initstate=0x0000000010007E6610C6402660301042 */ ;
    defparam mux_415_Mux_33.initval = 128'h0000000010007E6610C6402660301042;
    ROM128X1A mux_415_Mux_32 (.AD0(n25685), .AD1(n1359), .AD2(n1358), 
            .AD3(n1357), .AD4(n1356), .AD5(n1355), .AD6(n1354), .DO0(n725)) /* synthesis initstate=0x000000000000663C1046622438201042 */ ;
    defparam mux_415_Mux_32.initval = 128'h000000000000663C1046622438201042;
    FD1S3AY en_19 (.D(n5151), .CK(clk_c), .Q(en_c));   // g:/fpga/mxo2/system/project/system_top.v(45[10] 48[20])
    defparam en_19.GSR = "ENABLED";
    OB led_pad_5 (.I(rgb_led2_c), .O(led[5]));   // g:/fpga/mxo2/system/project/system_top.v(6[29:32])
    OB led_pad_6 (.I(rgb_led2_c), .O(led[6]));   // g:/fpga/mxo2/system/project/system_top.v(6[29:32])
    ROM128X1A mux_415_Mux_27 (.AD0(n25685), .AD1(n1359), .AD2(n1358), 
            .AD3(n1357), .AD4(n1356), .AD5(n1355), .AD6(n1354), .DO0(n864)) /* synthesis initstate=0x000000003800087E087C3E207C7E103C */ ;
    defparam mux_415_Mux_27.initval = 128'h000000003800087E087C3E207C7E103C;
    ROM128X1A mux_415_Mux_26 (.AD0(n25685), .AD1(n1359), .AD2(n1358), 
            .AD3(n1357), .AD4(n1356), .AD5(n1355), .AD6(n1354), .DO0(n865)) /* synthesis initstate=0x000000003C0018660846622066061064 */ ;
    defparam mux_415_Mux_26.initval = 128'h000000003C0018660846622066061064;
    ROM128X1A mux_415_Mux_25 (.AD0(n25685), .AD1(n1359), .AD2(n1358), 
            .AD3(n1357), .AD4(n1356), .AD5(n1355), .AD6(n1354), .DO0(n998)) /* synthesis initstate=0x0000000004003E3E7F103E303C3E183C */ ;
    defparam mux_415_Mux_25.initval = 128'h0000000004003E3E7F103E303C3E183C;
    ROM128X1A mux_415_Mux_24 (.AD0(n25685), .AD1(n1359), .AD2(n1358), 
            .AD3(n1357), .AD4(n1356), .AD5(n1355), .AD6(n1354), .DO0(n999)) /* synthesis initstate=0x0000000004001C1C7F103E201C1C181C */ ;
    defparam mux_415_Mux_24.initval = 128'h0000000004001C1C7F103E201C1C181C;
    BB one_wire_pad (.I(one_wire_N_501), .T(n5709), .B(one_wire), .O(one_wire_out));   // g:/fpga/mxo2/system/project/ds18b20z.v(48[1] 165[4])
    ROM128X1A mux_415_Mux_18 (.AD0(n25685), .AD1(n1359), .AD2(n1358), 
            .AD3(n1357), .AD4(n1356), .AD5(n1355), .AD6(n1354), .DO0(n1139)) /* synthesis initstate=0x0000000018006136103E3E2430201843 */ ;
    defparam mux_415_Mux_18.initval = 128'h0000000018006136103E3E2430201843;
    ROM128X1A mux_415_Mux_17 (.AD0(n25685), .AD1(n1359), .AD2(n1358), 
            .AD3(n1357), .AD4(n1356), .AD5(n1355), .AD6(n1354), .DO0(n1140)) /* synthesis initstate=0x000000002C00612230041E2C20201843 */ ;
    defparam mux_415_Mux_17.initval = 128'h000000002C00612230041E2C20201843;
    ROM128X1A mux_415_Mux_16 (.AD0(n25685), .AD1(n1359), .AD2(n1358), 
            .AD3(n1357), .AD4(n1356), .AD5(n1355), .AD6(n1354), .DO0(n1141)) /* synthesis initstate=0x00000000040061622004022860601A43 */ ;
    defparam mux_415_Mux_16.initval = 128'h00000000040061622004022860601A43;
    ROM128X1A mux_415_Mux_15 (.AD0(n25685), .AD1(n1359), .AD2(n1358), 
            .AD3(n1357), .AD4(n1356), .AD5(n1355), .AD6(n1354), .DO0(n1142)) /* synthesis initstate=0x0000000044186162200C022862601A62 */ ;
    defparam mux_415_Mux_15.initval = 128'h0000000044186162200C022862601A62;
    ROM128X1A mux_415_Mux_14 (.AD0(n25685), .AD1(n1359), .AD2(n1358), 
            .AD3(n1357), .AD4(n1356), .AD5(n1355), .AD6(n1354), .DO0(n1143)) /* synthesis initstate=0x00000000401863622008023862631E62 */ ;
    defparam mux_415_Mux_14.initval = 128'h00000000401863622008023862631E62;
    ROM128X1A mux_415_Mux_13 (.AD0(n25685), .AD1(n1359), .AD2(n1358), 
            .AD3(n1357), .AD4(n1356), .AD5(n1355), .AD6(n1354), .DO0(n1144)) /* synthesis initstate=0x00000000001863626008023062621C22 */ ;
    defparam mux_415_Mux_13.initval = 128'h00000000001863626008023062621C22;
    ROM128X1A mux_415_Mux_12 (.AD0(n25685), .AD1(n1359), .AD2(n1358), 
            .AD3(n1357), .AD4(n1356), .AD5(n1355), .AD6(n1354), .DO0(n1145)) /* synthesis initstate=0x00000000001836224018023026261826 */ ;
    defparam mux_415_Mux_12.initval = 128'h00000000001836224018023026261826;
    ROM128X1A mux_415_Mux_11 (.AD0(n25685), .AD1(n1359), .AD2(n1358), 
            .AD3(n1357), .AD4(n1356), .AD5(n1355), .AD6(n1354), .DO0(n1278)) /* synthesis initstate=0x000000002E1808630C42632062061822 */ ;
    defparam mux_415_Mux_11.initval = 128'h000000002E1808630C42632062061822;
    ROM128X1A mux_415_Mux_10 (.AD0(n25685), .AD1(n1359), .AD2(n1358), 
            .AD3(n1357), .AD4(n1356), .AD5(n1355), .AD6(n1354), .DO0(n1279)) /* synthesis initstate=0x000000002A1818430843617F63041862 */ ;
    defparam mux_415_Mux_10.initval = 128'h000000002A1818430843617F63041862;
    ROM128X1A mux_415_Mux_9 (.AD0(n25685), .AD1(n1359), .AD2(n1358), .AD3(n1357), 
            .AD4(n1356), .AD5(n1355), .AD6(n1354), .DO0(n1280)) /* synthesis initstate=0x000000004B1818410843607F420C1862 */ ;
    defparam mux_415_Mux_9.initval = 128'h000000004B1818410843607F420C1862;
    ROM128X1A mux_415_Mux_8 (.AD0(n25685), .AD1(n1359), .AD2(n1358), .AD3(n1357), 
            .AD4(n1356), .AD5(n1355), .AD6(n1354), .DO0(n1281)) /* synthesis initstate=0x00000000DB1810410843407F60081843 */ ;
    defparam mux_415_Mux_8.initval = 128'h00000000DB1810410843407F60081843;
    PFUMX i22155 (.BLUT(n25772), .ALUT(n25773), .C0(cnt_adj_5212[0]), 
          .Z(n25774));
    ROM128X1A mux_415_Mux_6 (.AD0(n25685), .AD1(n1359), .AD2(n1358), .AD3(n1357), 
            .AD4(n1356), .AD5(n1355), .AD6(n1354), .DO0(n1283)) /* synthesis initstate=0x0000000059003E631843602260101843 */ ;
    defparam mux_415_Mux_6.initval = 128'h0000000059003E631843602260101843;
    ROM128X1A mux_415_Mux_5 (.AD0(n25685), .AD1(n1359), .AD2(n1358), .AD3(n1357), 
            .AD4(n1356), .AD5(n1355), .AD6(n1354), .DO0(n1284)) /* synthesis initstate=0x0000000008003E361842602230101843 */ ;
    defparam mux_415_Mux_5.initval = 128'h0000000008003E361842602230101843;
    ROM128X1A mux_415_Mux_4 (.AD0(n25685), .AD1(n1359), .AD2(n1358), .AD3(n1357), 
            .AD4(n1356), .AD5(n1355), .AD6(n1354), .DO0(n1285)) /* synthesis initstate=0x000000000000333E1066232638301843 */ ;
    defparam mux_415_Mux_4.initval = 128'h000000000000333E1066232638301843;
    ROM128X1A mux_415_Mux_1 (.AD0(n25685), .AD1(n1359), .AD2(n1358), .AD3(n1357), 
            .AD4(n1356), .AD5(n1355), .AD6(n1354), .DO0(n1424)) /* synthesis initstate=0x000000001C000C3E043E3E203E7E183E */ ;
    defparam mux_415_Mux_1.initval = 128'h000000001C000C3E043E3E203E7E183E;
    OB rgb_led2_pad_2 (.I(rgb_led2_c), .O(rgb_led2[2]));   // g:/fpga/mxo2/system/project/system_top.v(8[29:37])
    OB rgb_led1_pad_0 (.I(rgb_led2_c), .O(rgb_led1[0]));   // g:/fpga/mxo2/system/project/system_top.v(7[29:37])
    OB rgb_led1_pad_1 (.I(rgb_led2_c), .O(rgb_led1[1]));   // g:/fpga/mxo2/system/project/system_top.v(7[29:37])
    OB rgb_led1_pad_2 (.I(rgb_led2_c), .O(rgb_led1[2]));   // g:/fpga/mxo2/system/project/system_top.v(7[29:37])
    OB led_pad_0 (.I(rgb_led2_c), .O(led[0]));   // g:/fpga/mxo2/system/project/system_top.v(6[29:32])
    OB led_pad_1 (.I(rgb_led2_c), .O(led[1]));   // g:/fpga/mxo2/system/project/system_top.v(6[29:32])
    OB led_pad_2 (.I(rgb_led2_c), .O(led[2]));   // g:/fpga/mxo2/system/project/system_top.v(6[29:32])
    OB led_pad_3 (.I(rgb_led2_c), .O(led[3]));   // g:/fpga/mxo2/system/project/system_top.v(6[29:32])
    OB led_pad_4 (.I(rgb_led2_c), .O(led[4]));   // g:/fpga/mxo2/system/project/system_top.v(6[29:32])
    OB rgb_led2_pad_1 (.I(rgb_led2_c), .O(rgb_led2[1]));   // g:/fpga/mxo2/system/project/system_top.v(8[29:37])
    LUT4 i21405_2_lut_rep_320_3_lut_4_lut (.A(clk_1mhz), .B(n25765), .C(state[0]), 
         .D(state_back_2__N_261[2]), .Z(clk_c_enable_1433)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam i21405_2_lut_rep_320_3_lut_4_lut.init = 16'h0004;
    LUT4 n24759_bdd_2_lut_3_lut (.A(clk_1mhz), .B(n25765), .C(n25857), 
         .Z(clk_c_enable_132)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam n24759_bdd_2_lut_3_lut.init = 16'h4040;
    LUT4 i2_3_lut_4_lut (.A(clk_1mhz), .B(n25765), .C(en_c), .D(data_out[2]), 
         .Z(n20945)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam i2_3_lut_4_lut.init = 16'h0040;
    LUT4 i1_2_lut_rep_325_3_lut (.A(clk_1mhz), .B(n25765), .C(state_back_2__N_261[2]), 
         .Z(n25607)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam i1_2_lut_rep_325_3_lut.init = 16'hfbfb;
    LUT4 i21409_2_lut_3_lut_4_lut (.A(clk_1mhz), .B(n25765), .C(state[1]), 
         .D(state_back_2__N_261[2]), .Z(clk_c_enable_1437)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam i21409_2_lut_3_lut_4_lut.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut (.A(clk_1mhz), .B(n25765), .C(n25484), .D(rst_n_c), 
         .Z(clk_c_enable_686)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 i1_2_lut_3_lut (.A(clk_1mhz), .B(n25765), .C(en_c), .Z(clk_c_enable_931)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam i1_2_lut_3_lut.init = 16'h4040;
    LUT4 i1_2_lut_rep_336_3_lut (.A(clk_1mhz), .B(n25765), .C(rst_n_c), 
         .Z(n25618)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam i1_2_lut_rep_336_3_lut.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_284 (.A(clk_1mhz), .B(n25765), .C(n25453), 
         .Z(clk_c_enable_1439)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam i1_2_lut_3_lut_adj_284.init = 16'h4040;
    LUT4 i20793_2_lut_3_lut_4_lut (.A(clk_1mhz), .B(n25765), .C(cnt_read[2]), 
         .D(rst_n_c), .Z(n23656)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam i20793_2_lut_3_lut_4_lut.init = 16'h4000;
    FD1S3AX led_i1 (.D(n26780), .CK(clk_c), .Q(rgb_led2_c));   // g:/fpga/mxo2/system/project/system_top.v(36[10] 40[8])
    defparam led_i1.GSR = "ENABLED";
    LUT4 i31_4_lut_4_lut (.A(cnt_adj_5212[0]), .B(cnt_adj_5212[1]), .C(cnt_adj_5212[4]), 
         .D(cnt_adj_5212[2]), .Z(n12)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A (B (C)+!B ((D)+!C)))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(87[20] 90[14])
    defparam i31_4_lut_4_lut.init = 16'h0494;
    LUT4 i2_4_lut (.A(n28), .B(n4), .C(state_back_2__N_261[2]), .D(n16602), 
         .Z(clk_c_enable_117)) /* synthesis lut_function=(A (B)+!A !((C+(D))+!B)) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(45[14:24])
    defparam i2_4_lut.init = 16'h888c;
    LUT4 i1_4_lut (.A(n50), .B(n25706), .C(n25742), .D(n16451), .Z(n4)) /* synthesis lut_function=(A (B+(C+!(D)))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(45[14:24])
    defparam i1_4_lut.init = 16'ha8aa;
    LUT4 i21089_4_lut_4_lut (.A(cnt_adj_5212[0]), .B(cnt_adj_5212[1]), .C(cnt_adj_5212[2]), 
         .D(cnt_adj_5212[3]), .Z(n23966)) /* synthesis lut_function=(A (D)+!A !(B (C+!(D))+!B !(C (D)+!C !(D)))) */ ;
    defparam i21089_4_lut_4_lut.init = 16'hbe01;
    LUT4 i2234_3_lut (.A(ready), .B(n26793), .C(n15), .Z(clk_c_enable_659)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i2234_3_lut.init = 16'hecec;
    LUT4 i1_2_lut_rep_424 (.A(state_back_2__N_261[2]), .B(state[0]), .Z(n25706)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_424.init = 16'heeee;
    LUT4 i1_3_lut_4_lut (.A(state_back_2__N_261[2]), .B(state[0]), .C(n25689), 
         .D(cnt_init[2]), .Z(num_delay_19__N_369[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C+!(D)))) */ ;
    defparam i1_3_lut_4_lut.init = 16'hf0f1;
    LUT4 i2233_2_lut (.A(ready), .B(n26793), .Z(clk_c_enable_1399)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2233_2_lut.init = 16'heeee;
    LUT4 mux_123_Mux_5_i31_then_4_lut (.A(cnt_adj_5212[3]), .B(cnt_adj_5212[4]), 
         .C(cnt_adj_5212[1]), .D(cnt_adj_5212[2]), .Z(n25773)) /* synthesis lut_function=(!(A (B+(C (D)+!C !(D)))+!A (B+(C (D))))) */ ;
    defparam mux_123_Mux_5_i31_then_4_lut.init = 16'h0331;
    LUT4 mux_123_Mux_5_i31_else_4_lut (.A(cnt_adj_5212[3]), .B(cnt_adj_5212[4]), 
         .C(cnt_adj_5212[1]), .D(cnt_adj_5212[2]), .Z(n25772)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)+!C !(D)))+!A (B+!(C (D)+!C !(D))))) */ ;
    defparam mux_123_Mux_5_i31_else_4_lut.init = 16'h1a21;
    GSR GSR_INST (.GSR(rst_n_c));
    LUT4 i32_3_lut_3_lut_4_lut (.A(cnt_adj_5212[1]), .B(cnt_adj_5212[2]), 
         .C(cnt_adj_5212[4]), .D(cnt_adj_5212[0]), .Z(n15_adj_5200)) /* synthesis lut_function=(!(A ((D)+!C)+!A !(B (C+(D))+!B !((D)+!C)))) */ ;
    defparam i32_3_lut_3_lut_4_lut.init = 16'h44f0;
    time_generator time_generator_inst (.time_data({time_data}), .clk_c(clk_c), 
            .flag(flag), .n26780(n26780), .en_c(en_c), .key_c_1(key_c_1), 
            .key_c_0(key_c_0), .key_c_2(key_c_2), .\data_out[1] (data_out[1]), 
            .\tamp_out_11__N_478[3] (tamp_out_11__N_478[3]), .\data_out[2] (data_out[2]), 
            .tamp_out_11__N_483(tamp_out_11__N_483), .\data_out[0] (data_out[0]), 
            .tamp_out_11__N_489(tamp_out_11__N_489), .\data_length_reg[0] (data_length_reg[0]), 
            .n15(n15_adj_5201), .n5151(n5151), .GND_net(GND_net), .tamp_out_11__N_495(tamp_out_11__N_495)) /* synthesis syn_module_defined=1 */ ;   // g:/fpga/mxo2/system/project/system_top.v(51[16] 58[2])
    LUT4 i21351_2_lut_rep_469 (.A(cnt_adj_5212[0]), .B(cnt_adj_5212[1]), 
         .Z(n25751)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i21351_2_lut_rep_469.init = 16'h1111;
    LUT4 i21148_3_lut_4_lut (.A(cnt_adj_5212[0]), .B(cnt_adj_5212[1]), .C(cnt_adj_5212[2]), 
         .D(cnt_adj_5212[3]), .Z(n23973)) /* synthesis lut_function=(!(A (B (C+!(D))+!B ((D)+!C))+!A (B (C)+!B !(C (D))))) */ ;
    defparam i21148_3_lut_4_lut.init = 16'h1c24;
    LUT4 m1_lut (.Z(n26780)) /* synthesis lut_function=1, syn_instantiated=1 */ ;
    defparam m1_lut.init = 16'hffff;
    LUT4 i21090_4_lut_4_lut_4_lut_4_lut (.A(cnt_adj_5212[0]), .B(cnt_adj_5212[3]), 
         .C(cnt_adj_5212[1]), .D(cnt_adj_5212[2]), .Z(n23967)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C (D))))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(87[20] 90[14])
    defparam i21090_4_lut_4_lut_4_lut_4_lut.init = 16'h1575;
    LUT4 i21095_4_lut_4_lut_4_lut (.A(cnt_adj_5212[0]), .B(cnt_adj_5212[1]), 
         .C(cnt_adj_5212[2]), .D(cnt_adj_5212[3]), .Z(n23972)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A !(B (D)+!B (C (D)+!C !(D))))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(87[20] 90[14])
    defparam i21095_4_lut_4_lut_4_lut.init = 16'h5421;
    OLED12832 OLED12832_inst (.clk_c(clk_c), .oled_csn_c(oled_csn_c), .n25808(n25808), 
            .n1358(n1358), .n1359(n1359), .n1138(n1138), .n1278(n1278), 
            .n998(n998), .n579(n579), .n719(n719), .n439(n439), .n578(n578), 
            .n718(n718), .n438(n438), .n1357(n1357), .n1356(n1356), 
            .n23966(n23966), .n23967(n23967), .cnt({Open_0, Open_1, 
            Open_2, Open_3, Open_4, Open_5, Open_6, Open_7, Open_8, 
            Open_9, Open_10, cnt_adj_5212[4:0]}), .n1141(n1141), .n1281(n1281), 
            .n1140(n1140), .n1280(n1280), .time_data({time_data}), .\tamp_data[1] (tamp_data[1]), 
            .n865(n865), .n582(n582), .n722(n722), .n581(n581), .n721(n721), 
            .n1139(n1139), .n1279(n1279), .n999(n999), .n583(n583), 
            .n723(n723), .n580(n580), .n720(n720), .n1142(n1142), .n1282(n1282), 
            .n1424(n1424), .n1144(n1144), .n1284(n1284), .n1143(n1143), 
            .n1283(n1283), .n584(n584), .n724(n724), .n1355(n1355), 
            .n25751(n25751), .n1354(n1354), .n23974(n23974), .n23971(n23971), 
            .n22685(n22685), .GND_net(GND_net), .n25774(n25774), .\tamp_data[3] (tamp_data[3]), 
            .n25685(n25685), .n863(n863), .n1423(n1423), .n1425(n1425), 
            .\tamp_data[0] (tamp_data[0]), .\tamp_data[8] (tamp_data[8]), 
            .\tamp_data[4] (tamp_data[4]), .\tamp_data[6] (tamp_data[6]), 
            .n864(n864), .oled_dat_c(oled_dat_c), .n25826(n25826), .oled_clk_c(oled_clk_c), 
            .oled_dcn_c(oled_dcn_c), .\tamp_data[7] (tamp_data[7]), .\tamp_data[9] (tamp_data[9]), 
            .\tamp_data[5] (tamp_data[5]), .oled_rst_c(oled_rst_c), .\tamp_data[2] (tamp_data[2]), 
            .n1145(n1145), .n585(n585), .n725(n725), .n1285(n1285)) /* synthesis syn_module_defined=1 */ ;   // g:/fpga/mxo2/system/project/system_top.v(70[11] 80[2])
    LUT4 i1_4_lut_adj_285 (.A(n50), .B(state_back_2__N_261[2]), .C(n28), 
         .D(n37), .Z(clk_c_enable_684)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))) */ ;
    defparam i1_4_lut_adj_285.init = 16'ha2a0;
    LUT4 i21093_4_lut_4_lut_4_lut (.A(cnt_adj_5212[0]), .B(cnt_adj_5212[1]), 
         .C(cnt_adj_5212[2]), .D(cnt_adj_5212[3]), .Z(n23970)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C (D)+!C !(D))+!B !(C+(D))))) */ ;
    defparam i21093_4_lut_4_lut_4_lut.init = 16'h1570;
    LUT4 i21092_3_lut_4_lut_4_lut (.A(cnt_adj_5212[0]), .B(cnt_adj_5212[2]), 
         .C(cnt_adj_5212[1]), .D(cnt_adj_5212[3]), .Z(n23969)) /* synthesis lut_function=(A (B ((D)+!C))+!A (B (C (D))+!B (C (D)+!C !(D)))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(87[20] 90[14])
    defparam i21092_3_lut_4_lut_4_lut.init = 16'hd809;
    LUT4 mux_123_Mux_6_i31_3_lut_then_4_lut (.A(cnt_adj_5212[4]), .B(cnt_adj_5212[0]), 
         .C(cnt_adj_5212[1]), .D(cnt_adj_5212[2]), .Z(n25807)) /* synthesis lut_function=(!(A (C+(D))+!A !(B (C (D))+!B !((D)+!C)))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(87[20] 90[14])
    defparam mux_123_Mux_6_i31_3_lut_then_4_lut.init = 16'h401a;
    LUT4 mux_123_Mux_6_i31_3_lut_else_4_lut (.A(cnt_adj_5212[4]), .B(cnt_adj_5212[0]), 
         .C(cnt_adj_5212[1]), .D(cnt_adj_5212[2]), .Z(n25806)) /* synthesis lut_function=(!(A (B)+!A ((C+!(D))+!B))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(87[20] 90[14])
    defparam mux_123_Mux_6_i31_3_lut_else_4_lut.init = 16'h2622;
    LUT4 i1_4_lut_adj_286 (.A(n50), .B(state_back_2__N_261[2]), .C(n28), 
         .D(n29), .Z(clk_c_enable_688)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))) */ ;
    defparam i1_4_lut_adj_286.init = 16'ha2a0;
    PFUMX i22190 (.BLUT(n25824), .ALUT(n25825), .C0(cnt_adj_5212[1]), 
          .Z(n25826));
    beeper_control piano_out_I_0 (.\data_buffer[538] (data_buffer[538]), .n26793(n26793), 
            .\data_buffer[539] (data_buffer[539]), .\data_buffer[540] (data_buffer[540]), 
            .\data_buffer[544] (data_buffer[544]), .\data_buffer[545] (data_buffer[545]), 
            .\data_buffer[546] (data_buffer[546]), .\data_buffer[547] (data_buffer[547]), 
            .\data_buffer[548] (data_buffer[548]), .\data_buffer[552] (data_buffer[552]), 
            .\data_buffer[553] (data_buffer[553]), .\data_buffer[554] (data_buffer[554]), 
            .\data_buffer[555] (data_buffer[555]), .\data_buffer[556] (data_buffer[556]), 
            .\data_buffer[560] (data_buffer[560]), .\data_buffer[561] (data_buffer[561]), 
            .\data_buffer[562] (data_buffer[562]), .\data_buffer[563] (data_buffer[563]), 
            .\data_buffer[564] (data_buffer[564]), .\data_buffer[568] (data_buffer[568]), 
            .\data_buffer[160] (data_buffer[160]), .\data_buffer[569] (data_buffer[569]), 
            .\data_buffer[570] (data_buffer[570]), .\data_buffer[571] (data_buffer[571]), 
            .clk_c(clk_c), .\data_buffer[572] (data_buffer[572]), .\data_buffer[576] (data_buffer[576]), 
            .\data_buffer[577] (data_buffer[577]), .\data_buffer[416] (data_buffer[416]), 
            .\data_buffer[578] (data_buffer[578]), .\data_buffer[579] (data_buffer[579]), 
            .\data_buffer[580] (data_buffer[580]), .\data_buffer[584] (data_buffer[584]), 
            .\data_buffer[585] (data_buffer[585]), .\data_buffer[586] (data_buffer[586]), 
            .\data_buffer[587] (data_buffer[587]), .\data_buffer[588] (data_buffer[588]), 
            .\data_buffer[592] (data_buffer[592]), .\data_buffer[593] (data_buffer[593]), 
            .\data_buffer[594] (data_buffer[594]), .\data_buffer[595] (data_buffer[595]), 
            .\data_buffer[596] (data_buffer[596]), .\data_buffer[600] (data_buffer[600]), 
            .\data_buffer[601] (data_buffer[601]), .\data_buffer[602] (data_buffer[602]), 
            .\data_buffer[603] (data_buffer[603]), .\data_buffer[604] (data_buffer[604]), 
            .\data_buffer[608] (data_buffer[608]), .\data_buffer[609] (data_buffer[609]), 
            .\data_buffer[610] (data_buffer[610]), .\data_buffer[611] (data_buffer[611]), 
            .\data_buffer[612] (data_buffer[612]), .\data_buffer[616] (data_buffer[616]), 
            .\data_buffer[617] (data_buffer[617]), .\data_buffer[618] (data_buffer[618]), 
            .\data_buffer[619] (data_buffer[619]), .\data_buffer[620] (data_buffer[620]), 
            .\data_buffer[624] (data_buffer[624]), .\data_buffer[625] (data_buffer[625]), 
            .\data_buffer[626] (data_buffer[626]), .\data_buffer[627] (data_buffer[627]), 
            .\data_buffer[628] (data_buffer[628]), .data_length_reg({Open_11, 
            Open_12, Open_13, Open_14, Open_15, Open_16, Open_17, 
            Open_18, Open_19, data_length_reg[0]}), .n15(n15_adj_5201), 
            .\data_buffer[632] (data_buffer[632]), .\data_buffer[633] (data_buffer[633]), 
            .\data_buffer[634] (data_buffer[634]), .\data_buffer[635] (data_buffer[635]), 
            .\data_buffer[636] (data_buffer[636]), .\data_buffer[640] (data_buffer[640]), 
            .\data_buffer[641] (data_buffer[641]), .\data_buffer[642] (data_buffer[642]), 
            .\data_buffer[643] (data_buffer[643]), .\data_buffer[644] (data_buffer[644]), 
            .\data_buffer[648] (data_buffer[648]), .\data_buffer[649] (data_buffer[649]), 
            .\data_buffer[650] (data_buffer[650]), .\data_buffer[651] (data_buffer[651]), 
            .\data_buffer[652] (data_buffer[652]), .\data_buffer[656] (data_buffer[656]), 
            .\data_buffer[657] (data_buffer[657]), .\data_buffer[658] (data_buffer[658]), 
            .\data_buffer[659] (data_buffer[659]), .\data_buffer[660] (data_buffer[660]), 
            .\data_buffer[664] (data_buffer[664]), .\data_buffer[665] (data_buffer[665]), 
            .\data_buffer[666] (data_buffer[666]), .\data_buffer[667] (data_buffer[667]), 
            .\data_buffer[668] (data_buffer[668]), .\data_buffer[672] (data_buffer[672]), 
            .\data_buffer[673] (data_buffer[673]), .\data_buffer[674] (data_buffer[674]), 
            .\data_buffer[675] (data_buffer[675]), .\data_buffer[676] (data_buffer[676]), 
            .\data_buffer[680] (data_buffer[680]), .\data_buffer[681] (data_buffer[681]), 
            .\data_buffer[682] (data_buffer[682]), .\data_buffer[683] (data_buffer[683]), 
            .\data_buffer[684] (data_buffer[684]), .\data_buffer[688] (data_buffer[688]), 
            .\data_buffer[689] (data_buffer[689]), .\data_buffer[690] (data_buffer[690]), 
            .\data_buffer[691] (data_buffer[691]), .\data_buffer[692] (data_buffer[692]), 
            .\data_buffer[696] (data_buffer[696]), .\data_buffer[697] (data_buffer[697]), 
            .\data_buffer[698] (data_buffer[698]), .\data_buffer[699] (data_buffer[699]), 
            .\data_buffer[700] (data_buffer[700]), .\data_buffer[704] (data_buffer[704]), 
            .\data_buffer[705] (data_buffer[705]), .\data_buffer[706] (data_buffer[706]), 
            .\data_buffer[707] (data_buffer[707]), .\data_buffer[708] (data_buffer[708]), 
            .\data_buffer[712] (data_buffer[712]), .\data_buffer[713] (data_buffer[713]), 
            .\data_buffer[714] (data_buffer[714]), .\data_buffer[715] (data_buffer[715]), 
            .\data_buffer[716] (data_buffer[716]), .\data_buffer[720] (data_buffer[720]), 
            .\data_buffer[161] (data_buffer[161]), .\data_buffer[721] (data_buffer[721]), 
            .\data_buffer[722] (data_buffer[722]), .\data_buffer[723] (data_buffer[723]), 
            .\data_buffer[724] (data_buffer[724]), .\data_buffer[728] (data_buffer[728]), 
            .\data_buffer[729] (data_buffer[729]), .\data_buffer[730] (data_buffer[730]), 
            .\data_buffer[731] (data_buffer[731]), .\data_buffer[732] (data_buffer[732]), 
            .\data_buffer[736] (data_buffer[736]), .\data_buffer[737] (data_buffer[737]), 
            .\data_buffer[162] (data_buffer[162]), .\data_buffer[738] (data_buffer[738]), 
            .\data_buffer[739] (data_buffer[739]), .\data_buffer[740] (data_buffer[740]), 
            .\data_buffer[744] (data_buffer[744]), .\data_buffer[163] (data_buffer[163]), 
            .\data_buffer[745] (data_buffer[745]), .\data_buffer[746] (data_buffer[746]), 
            .\data_buffer[747] (data_buffer[747]), .\data_buffer[748] (data_buffer[748]), 
            .\data_buffer[752] (data_buffer[752]), .\data_buffer[753] (data_buffer[753]), 
            .\data_buffer[754] (data_buffer[754]), .\data_buffer[755] (data_buffer[755]), 
            .\data_buffer[756] (data_buffer[756]), .\data_buffer[760] (data_buffer[760]), 
            .\data_buffer[761] (data_buffer[761]), .\data_buffer[762] (data_buffer[762]), 
            .\data_buffer[763] (data_buffer[763]), .\data_buffer[764] (data_buffer[764]), 
            .\data_buffer[768] (data_buffer[768]), .\data_buffer[769] (data_buffer[769]), 
            .\data_buffer[770] (data_buffer[770]), .\data_buffer[771] (data_buffer[771]), 
            .\data_buffer[772] (data_buffer[772]), .\data_buffer[776] (data_buffer[776]), 
            .\data_buffer[777] (data_buffer[777]), .\data_buffer[778] (data_buffer[778]), 
            .\data_buffer[779] (data_buffer[779]), .\data_buffer[780] (data_buffer[780]), 
            .\data_buffer[784] (data_buffer[784]), .\data_buffer[785] (data_buffer[785]), 
            .\data_buffer[786] (data_buffer[786]), .\data_buffer[787] (data_buffer[787]), 
            .\data_buffer[788] (data_buffer[788]), .\data_buffer[792] (data_buffer[792]), 
            .\data_buffer[793] (data_buffer[793]), .\data_buffer[794] (data_buffer[794]), 
            .\data_buffer[164] (data_buffer[164]), .\data_buffer[795] (data_buffer[795]), 
            .\data_buffer[796] (data_buffer[796]), .\data_buffer[800] (data_buffer[800]), 
            .\data_buffer[801] (data_buffer[801]), .\data_buffer[802] (data_buffer[802]), 
            .\data_buffer[803] (data_buffer[803]), .\data_buffer[804] (data_buffer[804]), 
            .\data_buffer[808] (data_buffer[808]), .\data_buffer[809] (data_buffer[809]), 
            .\data_buffer[810] (data_buffer[810]), .\data_buffer[811] (data_buffer[811]), 
            .\data_buffer[812] (data_buffer[812]), .\data_buffer[816] (data_buffer[816]), 
            .\data_buffer[817] (data_buffer[817]), .\data_buffer[818] (data_buffer[818]), 
            .\data_buffer[819] (data_buffer[819]), .\data_buffer[820] (data_buffer[820]), 
            .\data_buffer[824] (data_buffer[824]), .\data_buffer[825] (data_buffer[825]), 
            .\data_buffer[826] (data_buffer[826]), .\data_buffer[827] (data_buffer[827]), 
            .\data_buffer[828] (data_buffer[828]), .\data_buffer[832] (data_buffer[832]), 
            .\data_buffer[833] (data_buffer[833]), .\data_buffer[834] (data_buffer[834]), 
            .\data_buffer[835] (data_buffer[835]), .\data_buffer[836] (data_buffer[836]), 
            .\data_buffer[840] (data_buffer[840]), .\data_buffer[841] (data_buffer[841]), 
            .\data_buffer[842] (data_buffer[842]), .\data_buffer[843] (data_buffer[843]), 
            .\data_buffer[844] (data_buffer[844]), .\data_buffer[848] (data_buffer[848]), 
            .\data_buffer[849] (data_buffer[849]), .\data_buffer[850] (data_buffer[850]), 
            .\data_buffer[851] (data_buffer[851]), .\data_buffer[852] (data_buffer[852]), 
            .\data_buffer[856] (data_buffer[856]), .\data_buffer[857] (data_buffer[857]), 
            .\data_buffer[858] (data_buffer[858]), .\data_buffer[859] (data_buffer[859]), 
            .\data_buffer[860] (data_buffer[860]), .\data_buffer[864] (data_buffer[864]), 
            .\data_buffer[865] (data_buffer[865]), .\data_buffer[866] (data_buffer[866]), 
            .\data_buffer[867] (data_buffer[867]), .\data_buffer[868] (data_buffer[868]), 
            .\data_buffer[872] (data_buffer[872]), .\data_buffer[873] (data_buffer[873]), 
            .\data_buffer[874] (data_buffer[874]), .\data_buffer[875] (data_buffer[875]), 
            .\data_buffer[876] (data_buffer[876]), .\data_buffer[880] (data_buffer[880]), 
            .\data_buffer[881] (data_buffer[881]), .\data_buffer[882] (data_buffer[882]), 
            .\data_buffer[883] (data_buffer[883]), .\data_buffer[884] (data_buffer[884]), 
            .\data_buffer[888] (data_buffer[888]), .\data_buffer[889] (data_buffer[889]), 
            .\data_buffer[890] (data_buffer[890]), .\data_buffer[891] (data_buffer[891]), 
            .\data_buffer[892] (data_buffer[892]), .\data_buffer[386] (data_buffer[386]), 
            .\data_buffer[896] (data_buffer[896]), .\data_buffer[897] (data_buffer[897]), 
            .\data_buffer[898] (data_buffer[898]), .\data_buffer[899] (data_buffer[899]), 
            .\data_buffer[900] (data_buffer[900]), .\data_buffer[904] (data_buffer[904]), 
            .\data_buffer[905] (data_buffer[905]), .\data_buffer[906] (data_buffer[906]), 
            .\data_buffer[907] (data_buffer[907]), .\data_buffer[908] (data_buffer[908]), 
            .\data_buffer[912] (data_buffer[912]), .\data_buffer[913] (data_buffer[913]), 
            .\data_buffer[914] (data_buffer[914]), .\data_buffer[915] (data_buffer[915]), 
            .\data_buffer[916] (data_buffer[916]), .\data_buffer[920] (data_buffer[920]), 
            .\data_buffer[921] (data_buffer[921]), .\data_buffer[922] (data_buffer[922]), 
            .\data_buffer[923] (data_buffer[923]), .\data_buffer[924] (data_buffer[924]), 
            .\data_buffer[928] (data_buffer[928]), .\data_buffer[929] (data_buffer[929]), 
            .\data_buffer[930] (data_buffer[930]), .\data_buffer[931] (data_buffer[931]), 
            .\data_buffer[932] (data_buffer[932]), .\data_buffer[168] (data_buffer[168]), 
            .\data_buffer[936] (data_buffer[936]), .\data_buffer[937] (data_buffer[937]), 
            .\data_buffer[938] (data_buffer[938]), .\data_buffer[939] (data_buffer[939]), 
            .\data_buffer[940] (data_buffer[940]), .\data_buffer[944] (data_buffer[944]), 
            .\data_buffer[945] (data_buffer[945]), .\data_buffer[946] (data_buffer[946]), 
            .\data_buffer[947] (data_buffer[947]), .\data_buffer[948] (data_buffer[948]), 
            .\data_buffer[169] (data_buffer[169]), .\data_buffer[170] (data_buffer[170]), 
            .\data_buffer[171] (data_buffer[171]), .\data_buffer[0] (data_buffer[0]), 
            .\data_buffer[387] (data_buffer[387]), .\data_buffer[172] (data_buffer[172]), 
            .\data_buffer[176] (data_buffer[176]), .\data_buffer[177] (data_buffer[177]), 
            .\data_buffer[178] (data_buffer[178]), .\data_buffer[956] (data_buffer[956]), 
            .\data_buffer[179] (data_buffer[179]), .\data_buffer[1] (data_buffer[1]), 
            .\data_buffer[2] (data_buffer[2]), .\data_buffer[3] (data_buffer[3]), 
            .\data_buffer[4] (data_buffer[4]), .\data_buffer[8] (data_buffer[8]), 
            .\data_buffer[9] (data_buffer[9]), .\data_buffer[10] (data_buffer[10]), 
            .\data_buffer[11] (data_buffer[11]), .\data_buffer[12] (data_buffer[12]), 
            .\data_buffer[16] (data_buffer[16]), .\data_buffer[17] (data_buffer[17]), 
            .\data_buffer[18] (data_buffer[18]), .\data_buffer[19] (data_buffer[19]), 
            .\data_buffer[20] (data_buffer[20]), .\data_buffer[24] (data_buffer[24]), 
            .\data_buffer[25] (data_buffer[25]), .\data_buffer[26] (data_buffer[26]), 
            .\data_buffer[27] (data_buffer[27]), .\data_buffer[28] (data_buffer[28]), 
            .\data_buffer[32] (data_buffer[32]), .\data_buffer[33] (data_buffer[33]), 
            .\data_buffer[955] (data_buffer[955]), .\data_buffer[34] (data_buffer[34]), 
            .\data_buffer[35] (data_buffer[35]), .\data_buffer[36] (data_buffer[36]), 
            .\data_buffer[40] (data_buffer[40]), .\data_buffer[41] (data_buffer[41]), 
            .\data_buffer[42] (data_buffer[42]), .\data_buffer[43] (data_buffer[43]), 
            .\data_buffer[44] (data_buffer[44]), .\data_buffer[48] (data_buffer[48]), 
            .\data_buffer[49] (data_buffer[49]), .\data_buffer[50] (data_buffer[50]), 
            .\data_buffer[51] (data_buffer[51]), .\data_buffer[52] (data_buffer[52]), 
            .\data_buffer[56] (data_buffer[56]), .\data_buffer[57] (data_buffer[57]), 
            .\data_buffer[58] (data_buffer[58]), .\data_buffer[954] (data_buffer[954]), 
            .\data_buffer[59] (data_buffer[59]), .\data_buffer[60] (data_buffer[60]), 
            .\data_buffer[388] (data_buffer[388]), .\data_buffer[64] (data_buffer[64]), 
            .\data_buffer[953] (data_buffer[953]), .\data_buffer[952] (data_buffer[952]), 
            .\data_buffer[65] (data_buffer[65]), .\data_buffer[180] (data_buffer[180]), 
            .\data_buffer[66] (data_buffer[66]), .\data_buffer[67] (data_buffer[67]), 
            .\data_buffer[68] (data_buffer[68]), .\data_buffer[72] (data_buffer[72]), 
            .\data_buffer[73] (data_buffer[73]), .\data_buffer[74] (data_buffer[74]), 
            .\data_buffer[75] (data_buffer[75]), .\data_buffer[76] (data_buffer[76]), 
            .\data_buffer[80] (data_buffer[80]), .\data_buffer[81] (data_buffer[81]), 
            .\data_buffer[82] (data_buffer[82]), .\data_buffer[83] (data_buffer[83]), 
            .\data_buffer[84] (data_buffer[84]), .\data_buffer[88] (data_buffer[88]), 
            .\data_buffer[184] (data_buffer[184]), .\data_buffer[89] (data_buffer[89]), 
            .\data_buffer[90] (data_buffer[90]), .\data_buffer[185] (data_buffer[185]), 
            .\data_buffer[91] (data_buffer[91]), .\data_buffer[92] (data_buffer[92]), 
            .\data_buffer[96] (data_buffer[96]), .\data_buffer[97] (data_buffer[97]), 
            .\data_buffer[98] (data_buffer[98]), .\data_buffer[99] (data_buffer[99]), 
            .\data_buffer[100] (data_buffer[100]), .\data_buffer[186] (data_buffer[186]), 
            .\data_buffer[104] (data_buffer[104]), .\data_buffer[105] (data_buffer[105]), 
            .\data_buffer[106] (data_buffer[106]), .\data_buffer[107] (data_buffer[107]), 
            .\data_buffer[108] (data_buffer[108]), .\data_buffer[112] (data_buffer[112]), 
            .\data_buffer[113] (data_buffer[113]), .\data_buffer[114] (data_buffer[114]), 
            .\data_buffer[115] (data_buffer[115]), .\data_buffer[116] (data_buffer[116]), 
            .\data_buffer[120] (data_buffer[120]), .\data_buffer[121] (data_buffer[121]), 
            .\data_buffer[122] (data_buffer[122]), .\data_buffer[123] (data_buffer[123]), 
            .\data_buffer[124] (data_buffer[124]), .\data_buffer[128] (data_buffer[128]), 
            .\data_buffer[129] (data_buffer[129]), .\data_buffer[187] (data_buffer[187]), 
            .\data_buffer[130] (data_buffer[130]), .\data_buffer[131] (data_buffer[131]), 
            .\data_buffer[132] (data_buffer[132]), .\data_buffer[136] (data_buffer[136]), 
            .\data_buffer[137] (data_buffer[137]), .\data_buffer[138] (data_buffer[138]), 
            .\data_buffer[139] (data_buffer[139]), .\data_buffer[140] (data_buffer[140]), 
            .\data_buffer[144] (data_buffer[144]), .\data_buffer[145] (data_buffer[145]), 
            .\data_buffer[146] (data_buffer[146]), .\data_buffer[147] (data_buffer[147]), 
            .\data_buffer[148] (data_buffer[148]), .\data_buffer[152] (data_buffer[152]), 
            .\data_buffer[153] (data_buffer[153]), .\data_buffer[154] (data_buffer[154]), 
            .\data_buffer[155] (data_buffer[155]), .\data_buffer[156] (data_buffer[156]), 
            .\data_buffer[188] (data_buffer[188]), .\data_buffer[392] (data_buffer[392]), 
            .\data_buffer[393] (data_buffer[393]), .\data_buffer[394] (data_buffer[394]), 
            .\data_buffer[192] (data_buffer[192]), .\data_buffer[193] (data_buffer[193]), 
            .\data_buffer[194] (data_buffer[194]), .\data_buffer[195] (data_buffer[195]), 
            .\data_buffer[196] (data_buffer[196]), .\data_buffer[200] (data_buffer[200]), 
            .\data_buffer[395] (data_buffer[395]), .\data_buffer[396] (data_buffer[396]), 
            .\data_buffer[201] (data_buffer[201]), .\data_buffer[202] (data_buffer[202]), 
            .\data_buffer[203] (data_buffer[203]), .\data_buffer[204] (data_buffer[204]), 
            .\data_buffer[208] (data_buffer[208]), .\data_buffer[417] (data_buffer[417]), 
            .\data_buffer[418] (data_buffer[418]), .\data_buffer[419] (data_buffer[419]), 
            .\data_buffer[420] (data_buffer[420]), .\data_buffer[400] (data_buffer[400]), 
            .\data_buffer[401] (data_buffer[401]), .\data_buffer[209] (data_buffer[209]), 
            .\data_buffer[210] (data_buffer[210]), .\data_buffer[424] (data_buffer[424]), 
            .\data_buffer[211] (data_buffer[211]), .\data_buffer[425] (data_buffer[425]), 
            .\data_buffer[212] (data_buffer[212]), .\data_buffer[426] (data_buffer[426]), 
            .\data_buffer[402] (data_buffer[402]), .\data_buffer[427] (data_buffer[427]), 
            .\data_buffer[428] (data_buffer[428]), .\data_buffer[216] (data_buffer[216]), 
            .\data_buffer[217] (data_buffer[217]), .\data_buffer[218] (data_buffer[218]), 
            .\data_buffer[219] (data_buffer[219]), .\data_buffer[432] (data_buffer[432]), 
            .\data_buffer[433] (data_buffer[433]), .\data_buffer[220] (data_buffer[220]), 
            .\data_buffer[434] (data_buffer[434]), .\data_buffer[435] (data_buffer[435]), 
            .\data_buffer[436] (data_buffer[436]), .\data_buffer[440] (data_buffer[440]), 
            .\data_buffer[224] (data_buffer[224]), .\data_buffer[225] (data_buffer[225]), 
            .\data_buffer[441] (data_buffer[441]), .\data_buffer[403] (data_buffer[403]), 
            .\data_buffer[226] (data_buffer[226]), .\data_buffer[227] (data_buffer[227]), 
            .\data_buffer[228] (data_buffer[228]), .\data_buffer[232] (data_buffer[232]), 
            .\data_buffer[233] (data_buffer[233]), .\data_buffer[234] (data_buffer[234]), 
            .\data_buffer[442] (data_buffer[442]), .\data_buffer[443] (data_buffer[443]), 
            .\data_buffer[404] (data_buffer[404]), .\data_buffer[444] (data_buffer[444]), 
            .\data_buffer[235] (data_buffer[235]), .\data_buffer[236] (data_buffer[236]), 
            .\data_buffer[408] (data_buffer[408]), .\data_buffer[240] (data_buffer[240]), 
            .\data_buffer[409] (data_buffer[409]), .\data_buffer[241] (data_buffer[241]), 
            .\data_buffer[448] (data_buffer[448]), .\data_buffer[242] (data_buffer[242]), 
            .\data_buffer[449] (data_buffer[449]), .\data_buffer[450] (data_buffer[450]), 
            .\data_buffer[243] (data_buffer[243]), .\data_buffer[451] (data_buffer[451]), 
            .\data_buffer[244] (data_buffer[244]), .\data_buffer[248] (data_buffer[248]), 
            .\data_buffer[452] (data_buffer[452]), .\data_buffer[249] (data_buffer[249]), 
            .\data_buffer[250] (data_buffer[250]), .\data_buffer[251] (data_buffer[251]), 
            .\data_buffer[252] (data_buffer[252]), .\data_buffer[256] (data_buffer[256]), 
            .\data_buffer[257] (data_buffer[257]), .\data_buffer[258] (data_buffer[258]), 
            .\data_buffer[259] (data_buffer[259]), .\data_buffer[260] (data_buffer[260]), 
            .\data_buffer[264] (data_buffer[264]), .\data_buffer[265] (data_buffer[265]), 
            .\data_buffer[266] (data_buffer[266]), .\data_buffer[267] (data_buffer[267]), 
            .\data_buffer[268] (data_buffer[268]), .\data_buffer[272] (data_buffer[272]), 
            .\data_buffer[456] (data_buffer[456]), .\data_buffer[273] (data_buffer[273]), 
            .\data_buffer[274] (data_buffer[274]), .\data_buffer[457] (data_buffer[457]), 
            .\data_buffer[275] (data_buffer[275]), .\data_buffer[276] (data_buffer[276]), 
            .\data_buffer[458] (data_buffer[458]), .data_length({data_length}), 
            .GND_net(GND_net), .\data_buffer[280] (data_buffer[280]), .\data_buffer[459] (data_buffer[459]), 
            .\data_buffer[460] (data_buffer[460]), .\data_buffer[281] (data_buffer[281]), 
            .\data_buffer[282] (data_buffer[282]), .\data_buffer[283] (data_buffer[283]), 
            .\data_buffer[284] (data_buffer[284]), .\data_buffer[288] (data_buffer[288]), 
            .\data_buffer[464] (data_buffer[464]), .\data_buffer[289] (data_buffer[289]), 
            .\data_buffer[465] (data_buffer[465]), .\data_buffer[290] (data_buffer[290]), 
            .\data_buffer[466] (data_buffer[466]), .\data_buffer[291] (data_buffer[291]), 
            .\data_buffer[292] (data_buffer[292]), .\data_buffer[296] (data_buffer[296]), 
            .\data_buffer[467] (data_buffer[467]), .\data_buffer[297] (data_buffer[297]), 
            .\data_buffer[298] (data_buffer[298]), .\data_buffer[468] (data_buffer[468]), 
            .\data_buffer[472] (data_buffer[472]), .\data_buffer[299] (data_buffer[299]), 
            .\data_buffer[300] (data_buffer[300]), .\data_buffer[304] (data_buffer[304]), 
            .\data_buffer[305] (data_buffer[305]), .\data_buffer[306] (data_buffer[306]), 
            .\data_buffer[307] (data_buffer[307]), .\data_buffer[308] (data_buffer[308]), 
            .\data_buffer[312] (data_buffer[312]), .\data_buffer[473] (data_buffer[473]), 
            .\data_buffer[313] (data_buffer[313]), .\data_buffer[314] (data_buffer[314]), 
            .\data_buffer[315] (data_buffer[315]), .\data_buffer[474] (data_buffer[474]), 
            .\data_buffer[316] (data_buffer[316]), .\data_buffer[475] (data_buffer[475]), 
            .\data_buffer[320] (data_buffer[320]), .\data_buffer[321] (data_buffer[321]), 
            .\data_buffer[476] (data_buffer[476]), .\data_buffer[480] (data_buffer[480]), 
            .\data_buffer[322] (data_buffer[322]), .\data_buffer[323] (data_buffer[323]), 
            .\data_buffer[324] (data_buffer[324]), .\data_buffer[481] (data_buffer[481]), 
            .\data_buffer[328] (data_buffer[328]), .\data_buffer[329] (data_buffer[329]), 
            .\data_buffer[330] (data_buffer[330]), .\data_buffer[331] (data_buffer[331]), 
            .\data_buffer[482] (data_buffer[482]), .\data_buffer[483] (data_buffer[483]), 
            .\data_buffer[484] (data_buffer[484]), .\data_buffer[332] (data_buffer[332]), 
            .\data_buffer[488] (data_buffer[488]), .\data_buffer[336] (data_buffer[336]), 
            .\data_buffer[337] (data_buffer[337]), .\data_buffer[489] (data_buffer[489]), 
            .\data_buffer[338] (data_buffer[338]), .\data_buffer[490] (data_buffer[490]), 
            .\data_buffer[339] (data_buffer[339]), .\data_buffer[491] (data_buffer[491]), 
            .\data_buffer[340] (data_buffer[340]), .\data_buffer[344] (data_buffer[344]), 
            .\data_buffer[492] (data_buffer[492]), .\data_buffer[345] (data_buffer[345]), 
            .\data_buffer[496] (data_buffer[496]), .\data_buffer[497] (data_buffer[497]), 
            .\data_buffer[346] (data_buffer[346]), .\data_buffer[347] (data_buffer[347]), 
            .\data_buffer[498] (data_buffer[498]), .\data_buffer[499] (data_buffer[499]), 
            .\data_buffer[500] (data_buffer[500]), .\data_buffer[348] (data_buffer[348]), 
            .\data_buffer[352] (data_buffer[352]), .\data_buffer[353] (data_buffer[353]), 
            .\data_buffer[354] (data_buffer[354]), .\data_buffer[355] (data_buffer[355]), 
            .\data_buffer[356] (data_buffer[356]), .\data_buffer[504] (data_buffer[504]), 
            .\data_buffer[360] (data_buffer[360]), .\data_buffer[361] (data_buffer[361]), 
            .\data_buffer[505] (data_buffer[505]), .\data_buffer[506] (data_buffer[506]), 
            .\data_buffer[362] (data_buffer[362]), .\data_buffer[507] (data_buffer[507]), 
            .\data_buffer[363] (data_buffer[363]), .\data_buffer[508] (data_buffer[508]), 
            .\data_buffer[364] (data_buffer[364]), .\data_buffer[368] (data_buffer[368]), 
            .\data_buffer[369] (data_buffer[369]), .\data_buffer[512] (data_buffer[512]), 
            .\data_buffer[513] (data_buffer[513]), .\data_buffer[514] (data_buffer[514]), 
            .\data_buffer[515] (data_buffer[515]), .\data_buffer[370] (data_buffer[370]), 
            .\data_buffer[516] (data_buffer[516]), .\data_buffer[520] (data_buffer[520]), 
            .\data_buffer[371] (data_buffer[371]), .\data_buffer[521] (data_buffer[521]), 
            .\data_buffer[372] (data_buffer[372]), .\data_buffer[522] (data_buffer[522]), 
            .\data_buffer[523] (data_buffer[523]), .\data_buffer[524] (data_buffer[524]), 
            .\data_buffer[376] (data_buffer[376]), .\data_buffer[528] (data_buffer[528]), 
            .\data_buffer[529] (data_buffer[529]), .\data_buffer[530] (data_buffer[530]), 
            .\data_buffer[531] (data_buffer[531]), .\data_buffer[532] (data_buffer[532]), 
            .\data_buffer[536] (data_buffer[536]), .\data_buffer[537] (data_buffer[537]), 
            .\data_buffer[377] (data_buffer[377]), .\data_buffer[378] (data_buffer[378]), 
            .\data_buffer[379] (data_buffer[379]), .\data_buffer[380] (data_buffer[380]), 
            .\data_buffer[410] (data_buffer[410]), .\data_buffer[411] (data_buffer[411]), 
            .\data_buffer[412] (data_buffer[412]), .\data_buffer[384] (data_buffer[384]), 
            .\data_buffer[385] (data_buffer[385]), .piano_out_c(piano_out_c)) /* synthesis syn_module_defined=1 */ ;   // g:/fpga/mxo2/system/project/system_top.v(104[16] 113[2])
    uart_top uart_top_inst (.\data_buffer[432] (data_buffer[432]), .clk_c(clk_c), 
            .clk_c_enable_659(clk_c_enable_659), .\data_buffer[424] (data_buffer[424]), 
            .\data_buffer[0] (data_buffer[0]), .\data_buffer[956] (data_buffer[956]), 
            .\data_buffer[948] (data_buffer[948]), .\data_buffer[955] (data_buffer[955]), 
            .\data_buffer[947] (data_buffer[947]), .\data_buffer[954] (data_buffer[954]), 
            .\data_buffer[946] (data_buffer[946]), .\data_buffer[953] (data_buffer[953]), 
            .\data_buffer[945] (data_buffer[945]), .\data_buffer[952] (data_buffer[952]), 
            .\data_buffer[944] (data_buffer[944]), .\data_buffer[940] (data_buffer[940]), 
            .\data_buffer[939] (data_buffer[939]), .\data_buffer[938] (data_buffer[938]), 
            .\data_buffer[937] (data_buffer[937]), .\data_buffer[936] (data_buffer[936]), 
            .\data_buffer[932] (data_buffer[932]), .\data_buffer[931] (data_buffer[931]), 
            .\data_buffer[930] (data_buffer[930]), .\data_buffer[929] (data_buffer[929]), 
            .\data_buffer[928] (data_buffer[928]), .\data_buffer[924] (data_buffer[924]), 
            .\data_buffer[923] (data_buffer[923]), .\data_buffer[922] (data_buffer[922]), 
            .\data_buffer[921] (data_buffer[921]), .\data_buffer[920] (data_buffer[920]), 
            .\data_buffer[916] (data_buffer[916]), .\data_buffer[915] (data_buffer[915]), 
            .\data_buffer[914] (data_buffer[914]), .\data_buffer[913] (data_buffer[913]), 
            .\data_buffer[912] (data_buffer[912]), .\data_buffer[908] (data_buffer[908]), 
            .\data_buffer[907] (data_buffer[907]), .\data_buffer[906] (data_buffer[906]), 
            .\data_buffer[905] (data_buffer[905]), .\data_buffer[904] (data_buffer[904]), 
            .\data_buffer[900] (data_buffer[900]), .\data_buffer[899] (data_buffer[899]), 
            .\data_buffer[898] (data_buffer[898]), .\data_buffer[897] (data_buffer[897]), 
            .\data_buffer[896] (data_buffer[896]), .\data_buffer[892] (data_buffer[892]), 
            .\data_buffer[891] (data_buffer[891]), .\data_buffer[428] (data_buffer[428]), 
            .\data_buffer[420] (data_buffer[420]), .\data_buffer[427] (data_buffer[427]), 
            .\data_buffer[419] (data_buffer[419]), .\data_buffer[890] (data_buffer[890]), 
            .\data_buffer[889] (data_buffer[889]), .\data_buffer[888] (data_buffer[888]), 
            .\data_buffer[884] (data_buffer[884]), .\data_buffer[883] (data_buffer[883]), 
            .\data_buffer[882] (data_buffer[882]), .\data_buffer[881] (data_buffer[881]), 
            .\data_buffer[880] (data_buffer[880]), .\data_buffer[876] (data_buffer[876]), 
            .\data_buffer[875] (data_buffer[875]), .\data_buffer[874] (data_buffer[874]), 
            .\data_buffer[873] (data_buffer[873]), .\data_buffer[872] (data_buffer[872]), 
            .\data_buffer[868] (data_buffer[868]), .\data_buffer[867] (data_buffer[867]), 
            .\data_buffer[866] (data_buffer[866]), .\data_buffer[865] (data_buffer[865]), 
            .\data_buffer[864] (data_buffer[864]), .\data_buffer[860] (data_buffer[860]), 
            .\data_buffer[859] (data_buffer[859]), .\data_buffer[858] (data_buffer[858]), 
            .\data_buffer[857] (data_buffer[857]), .\data_buffer[856] (data_buffer[856]), 
            .\data_buffer[852] (data_buffer[852]), .\data_buffer[851] (data_buffer[851]), 
            .\data_buffer[850] (data_buffer[850]), .\data_buffer[849] (data_buffer[849]), 
            .\data_buffer[848] (data_buffer[848]), .\data_buffer[844] (data_buffer[844]), 
            .\data_buffer[843] (data_buffer[843]), .\data_buffer[842] (data_buffer[842]), 
            .\data_buffer[841] (data_buffer[841]), .\data_buffer[840] (data_buffer[840]), 
            .\data_buffer[836] (data_buffer[836]), .\data_buffer[835] (data_buffer[835]), 
            .\data_buffer[834] (data_buffer[834]), .\data_buffer[833] (data_buffer[833]), 
            .\data_buffer[832] (data_buffer[832]), .\data_buffer[828] (data_buffer[828]), 
            .\data_buffer[827] (data_buffer[827]), .\data_buffer[826] (data_buffer[826]), 
            .\data_buffer[825] (data_buffer[825]), .\data_buffer[824] (data_buffer[824]), 
            .\data_buffer[820] (data_buffer[820]), .\data_buffer[819] (data_buffer[819]), 
            .\data_buffer[818] (data_buffer[818]), .\data_buffer[817] (data_buffer[817]), 
            .\data_buffer[816] (data_buffer[816]), .\data_buffer[812] (data_buffer[812]), 
            .\data_buffer[811] (data_buffer[811]), .\data_buffer[810] (data_buffer[810]), 
            .\data_buffer[809] (data_buffer[809]), .\data_buffer[808] (data_buffer[808]), 
            .\data_buffer[804] (data_buffer[804]), .\data_buffer[803] (data_buffer[803]), 
            .\data_buffer[802] (data_buffer[802]), .\data_buffer[801] (data_buffer[801]), 
            .\data_buffer[800] (data_buffer[800]), .\data_buffer[796] (data_buffer[796]), 
            .\data_buffer[795] (data_buffer[795]), .\data_buffer[794] (data_buffer[794]), 
            .\data_buffer[793] (data_buffer[793]), .\data_buffer[792] (data_buffer[792]), 
            .n26780(n26780), .\data_buffer[788] (data_buffer[788]), .\data_buffer[787] (data_buffer[787]), 
            .\data_buffer[786] (data_buffer[786]), .\data_buffer[785] (data_buffer[785]), 
            .\data_buffer[784] (data_buffer[784]), .\data_buffer[780] (data_buffer[780]), 
            .\data_buffer[779] (data_buffer[779]), .\data_buffer[778] (data_buffer[778]), 
            .\data_buffer[777] (data_buffer[777]), .\data_buffer[776] (data_buffer[776]), 
            .\data_buffer[772] (data_buffer[772]), .\data_buffer[771] (data_buffer[771]), 
            .\data_buffer[770] (data_buffer[770]), .\data_buffer[769] (data_buffer[769]), 
            .\data_buffer[768] (data_buffer[768]), .\data_buffer[764] (data_buffer[764]), 
            .\data_buffer[763] (data_buffer[763]), .\data_buffer[762] (data_buffer[762]), 
            .\data_buffer[761] (data_buffer[761]), .\data_buffer[760] (data_buffer[760]), 
            .\data_buffer[756] (data_buffer[756]), .\data_buffer[755] (data_buffer[755]), 
            .\data_buffer[754] (data_buffer[754]), .\data_buffer[753] (data_buffer[753]), 
            .\data_buffer[752] (data_buffer[752]), .\data_buffer[748] (data_buffer[748]), 
            .\data_buffer[747] (data_buffer[747]), .\data_buffer[746] (data_buffer[746]), 
            .\data_buffer[745] (data_buffer[745]), .\data_buffer[744] (data_buffer[744]), 
            .\data_buffer[740] (data_buffer[740]), .\data_buffer[739] (data_buffer[739]), 
            .\data_buffer[738] (data_buffer[738]), .\data_buffer[737] (data_buffer[737]), 
            .\data_buffer[736] (data_buffer[736]), .\data_buffer[732] (data_buffer[732]), 
            .\data_buffer[731] (data_buffer[731]), .\data_buffer[730] (data_buffer[730]), 
            .\data_buffer[729] (data_buffer[729]), .\data_buffer[728] (data_buffer[728]), 
            .\data_buffer[724] (data_buffer[724]), .\data_buffer[723] (data_buffer[723]), 
            .\data_buffer[722] (data_buffer[722]), .\data_buffer[721] (data_buffer[721]), 
            .\data_buffer[720] (data_buffer[720]), .\data_buffer[716] (data_buffer[716]), 
            .\data_buffer[715] (data_buffer[715]), .\data_buffer[714] (data_buffer[714]), 
            .\data_buffer[713] (data_buffer[713]), .\data_buffer[712] (data_buffer[712]), 
            .\data_buffer[708] (data_buffer[708]), .\data_buffer[707] (data_buffer[707]), 
            .\data_buffer[706] (data_buffer[706]), .\data_buffer[705] (data_buffer[705]), 
            .\data_buffer[704] (data_buffer[704]), .\data_buffer[700] (data_buffer[700]), 
            .\data_buffer[699] (data_buffer[699]), .\data_buffer[698] (data_buffer[698]), 
            .\data_buffer[697] (data_buffer[697]), .\data_buffer[696] (data_buffer[696]), 
            .\data_buffer[692] (data_buffer[692]), .\data_buffer[691] (data_buffer[691]), 
            .\data_buffer[690] (data_buffer[690]), .\data_buffer[689] (data_buffer[689]), 
            .\data_buffer[688] (data_buffer[688]), .\data_buffer[684] (data_buffer[684]), 
            .\data_buffer[683] (data_buffer[683]), .\data_buffer[682] (data_buffer[682]), 
            .\data_buffer[681] (data_buffer[681]), .\data_buffer[680] (data_buffer[680]), 
            .\data_buffer[676] (data_buffer[676]), .\data_buffer[675] (data_buffer[675]), 
            .\data_buffer[674] (data_buffer[674]), .\data_buffer[673] (data_buffer[673]), 
            .\data_buffer[672] (data_buffer[672]), .\data_buffer[668] (data_buffer[668]), 
            .\data_buffer[667] (data_buffer[667]), .\data_buffer[666] (data_buffer[666]), 
            .\data_buffer[665] (data_buffer[665]), .\data_buffer[664] (data_buffer[664]), 
            .\data_buffer[660] (data_buffer[660]), .\data_buffer[659] (data_buffer[659]), 
            .\data_buffer[658] (data_buffer[658]), .\data_buffer[657] (data_buffer[657]), 
            .\data_buffer[656] (data_buffer[656]), .\data_buffer[652] (data_buffer[652]), 
            .\data_buffer[651] (data_buffer[651]), .\data_buffer[650] (data_buffer[650]), 
            .\data_buffer[649] (data_buffer[649]), .\data_buffer[648] (data_buffer[648]), 
            .\data_buffer[644] (data_buffer[644]), .\data_buffer[643] (data_buffer[643]), 
            .\data_buffer[642] (data_buffer[642]), .\data_buffer[641] (data_buffer[641]), 
            .\data_buffer[640] (data_buffer[640]), .\data_buffer[636] (data_buffer[636]), 
            .\data_buffer[635] (data_buffer[635]), .\data_buffer[634] (data_buffer[634]), 
            .\data_buffer[633] (data_buffer[633]), .\data_buffer[632] (data_buffer[632]), 
            .\data_buffer[628] (data_buffer[628]), .\data_buffer[627] (data_buffer[627]), 
            .\data_buffer[626] (data_buffer[626]), .\data_buffer[625] (data_buffer[625]), 
            .\data_buffer[624] (data_buffer[624]), .\data_buffer[620] (data_buffer[620]), 
            .\data_buffer[619] (data_buffer[619]), .\data_buffer[618] (data_buffer[618]), 
            .\data_buffer[617] (data_buffer[617]), .\data_buffer[616] (data_buffer[616]), 
            .\data_buffer[612] (data_buffer[612]), .\data_buffer[611] (data_buffer[611]), 
            .\data_buffer[610] (data_buffer[610]), .\data_buffer[609] (data_buffer[609]), 
            .\data_buffer[608] (data_buffer[608]), .\data_buffer[604] (data_buffer[604]), 
            .\data_buffer[603] (data_buffer[603]), .\data_buffer[602] (data_buffer[602]), 
            .\data_buffer[601] (data_buffer[601]), .\data_buffer[600] (data_buffer[600]), 
            .\data_buffer[596] (data_buffer[596]), .\data_buffer[595] (data_buffer[595]), 
            .\data_buffer[594] (data_buffer[594]), .\data_buffer[593] (data_buffer[593]), 
            .\data_buffer[592] (data_buffer[592]), .\data_buffer[588] (data_buffer[588]), 
            .\data_buffer[587] (data_buffer[587]), .\data_buffer[586] (data_buffer[586]), 
            .\data_buffer[585] (data_buffer[585]), .\data_buffer[584] (data_buffer[584]), 
            .\data_buffer[580] (data_buffer[580]), .\data_buffer[579] (data_buffer[579]), 
            .\data_buffer[578] (data_buffer[578]), .\data_buffer[577] (data_buffer[577]), 
            .\data_buffer[576] (data_buffer[576]), .\data_buffer[572] (data_buffer[572]), 
            .\data_buffer[571] (data_buffer[571]), .\data_buffer[570] (data_buffer[570]), 
            .\data_buffer[569] (data_buffer[569]), .\data_buffer[568] (data_buffer[568]), 
            .\data_buffer[564] (data_buffer[564]), .\data_buffer[563] (data_buffer[563]), 
            .\data_buffer[562] (data_buffer[562]), .\data_buffer[561] (data_buffer[561]), 
            .\data_buffer[560] (data_buffer[560]), .\data_buffer[556] (data_buffer[556]), 
            .\data_buffer[555] (data_buffer[555]), .\data_buffer[554] (data_buffer[554]), 
            .\data_buffer[553] (data_buffer[553]), .\data_buffer[552] (data_buffer[552]), 
            .\data_buffer[548] (data_buffer[548]), .\data_buffer[547] (data_buffer[547]), 
            .\data_buffer[546] (data_buffer[546]), .\data_buffer[545] (data_buffer[545]), 
            .\data_buffer[544] (data_buffer[544]), .\data_buffer[540] (data_buffer[540]), 
            .\data_buffer[539] (data_buffer[539]), .\data_buffer[538] (data_buffer[538]), 
            .\data_buffer[537] (data_buffer[537]), .\data_buffer[536] (data_buffer[536]), 
            .\data_buffer[532] (data_buffer[532]), .\data_buffer[531] (data_buffer[531]), 
            .\data_buffer[530] (data_buffer[530]), .\data_buffer[529] (data_buffer[529]), 
            .\data_buffer[528] (data_buffer[528]), .\data_buffer[524] (data_buffer[524]), 
            .\data_buffer[523] (data_buffer[523]), .\data_buffer[522] (data_buffer[522]), 
            .\data_buffer[521] (data_buffer[521]), .\data_buffer[520] (data_buffer[520]), 
            .\data_buffer[516] (data_buffer[516]), .\data_buffer[515] (data_buffer[515]), 
            .\data_buffer[514] (data_buffer[514]), .\data_buffer[513] (data_buffer[513]), 
            .\data_buffer[512] (data_buffer[512]), .\data_buffer[508] (data_buffer[508]), 
            .\data_buffer[507] (data_buffer[507]), .\data_buffer[506] (data_buffer[506]), 
            .\data_buffer[505] (data_buffer[505]), .\data_buffer[504] (data_buffer[504]), 
            .\data_buffer[500] (data_buffer[500]), .\data_buffer[499] (data_buffer[499]), 
            .\data_buffer[498] (data_buffer[498]), .\data_buffer[497] (data_buffer[497]), 
            .\data_buffer[496] (data_buffer[496]), .\data_buffer[492] (data_buffer[492]), 
            .\data_buffer[491] (data_buffer[491]), .\data_buffer[490] (data_buffer[490]), 
            .\data_buffer[489] (data_buffer[489]), .\data_buffer[488] (data_buffer[488]), 
            .\data_buffer[484] (data_buffer[484]), .\data_buffer[483] (data_buffer[483]), 
            .\data_buffer[482] (data_buffer[482]), .\data_buffer[481] (data_buffer[481]), 
            .\data_buffer[480] (data_buffer[480]), .\data_buffer[476] (data_buffer[476]), 
            .\data_buffer[475] (data_buffer[475]), .\data_buffer[474] (data_buffer[474]), 
            .\data_buffer[473] (data_buffer[473]), .\data_buffer[472] (data_buffer[472]), 
            .\data_buffer[468] (data_buffer[468]), .\data_buffer[467] (data_buffer[467]), 
            .\data_buffer[466] (data_buffer[466]), .\data_buffer[465] (data_buffer[465]), 
            .\data_buffer[464] (data_buffer[464]), .\data_buffer[460] (data_buffer[460]), 
            .\data_buffer[459] (data_buffer[459]), .\data_buffer[458] (data_buffer[458]), 
            .\data_buffer[457] (data_buffer[457]), .\data_buffer[456] (data_buffer[456]), 
            .\data_buffer[452] (data_buffer[452]), .\data_buffer[451] (data_buffer[451]), 
            .\data_buffer[450] (data_buffer[450]), .\data_buffer[449] (data_buffer[449]), 
            .\data_buffer[448] (data_buffer[448]), .\data_buffer[444] (data_buffer[444]), 
            .\data_buffer[443] (data_buffer[443]), .\data_buffer[442] (data_buffer[442]), 
            .\data_buffer[441] (data_buffer[441]), .\data_buffer[440] (data_buffer[440]), 
            .\data_buffer[436] (data_buffer[436]), .\data_buffer[435] (data_buffer[435]), 
            .\data_buffer[434] (data_buffer[434]), .\data_buffer[433] (data_buffer[433]), 
            .\data_buffer[426] (data_buffer[426]), .\data_buffer[425] (data_buffer[425]), 
            .\data_buffer[418] (data_buffer[418]), .\data_buffer[417] (data_buffer[417]), 
            .\data_buffer[416] (data_buffer[416]), .\data_buffer[412] (data_buffer[412]), 
            .\data_buffer[411] (data_buffer[411]), .\data_buffer[410] (data_buffer[410]), 
            .\data_buffer[409] (data_buffer[409]), .\data_buffer[408] (data_buffer[408]), 
            .\data_buffer[404] (data_buffer[404]), .\data_buffer[403] (data_buffer[403]), 
            .\data_buffer[402] (data_buffer[402]), .\data_buffer[401] (data_buffer[401]), 
            .\data_buffer[400] (data_buffer[400]), .\data_buffer[396] (data_buffer[396]), 
            .\data_buffer[395] (data_buffer[395]), .\data_buffer[394] (data_buffer[394]), 
            .\data_buffer[393] (data_buffer[393]), .\data_buffer[392] (data_buffer[392]), 
            .\data_buffer[388] (data_buffer[388]), .\data_buffer[387] (data_buffer[387]), 
            .\data_buffer[386] (data_buffer[386]), .\data_buffer[385] (data_buffer[385]), 
            .\data_buffer[384] (data_buffer[384]), .\data_buffer[380] (data_buffer[380]), 
            .\data_buffer[379] (data_buffer[379]), .\data_buffer[378] (data_buffer[378]), 
            .\data_buffer[377] (data_buffer[377]), .\data_buffer[376] (data_buffer[376]), 
            .\data_buffer[372] (data_buffer[372]), .\data_buffer[371] (data_buffer[371]), 
            .\data_buffer[370] (data_buffer[370]), .\data_buffer[369] (data_buffer[369]), 
            .\data_buffer[368] (data_buffer[368]), .\data_buffer[364] (data_buffer[364]), 
            .\data_buffer[363] (data_buffer[363]), .\data_buffer[362] (data_buffer[362]), 
            .\data_buffer[361] (data_buffer[361]), .\data_buffer[360] (data_buffer[360]), 
            .\data_buffer[356] (data_buffer[356]), .\data_buffer[355] (data_buffer[355]), 
            .\data_buffer[354] (data_buffer[354]), .\data_buffer[353] (data_buffer[353]), 
            .\data_buffer[352] (data_buffer[352]), .\data_buffer[348] (data_buffer[348]), 
            .\data_buffer[347] (data_buffer[347]), .\data_buffer[346] (data_buffer[346]), 
            .\data_buffer[345] (data_buffer[345]), .\data_buffer[344] (data_buffer[344]), 
            .\data_buffer[340] (data_buffer[340]), .\data_buffer[339] (data_buffer[339]), 
            .\data_buffer[338] (data_buffer[338]), .\data_buffer[337] (data_buffer[337]), 
            .\data_buffer[336] (data_buffer[336]), .\data_buffer[332] (data_buffer[332]), 
            .\data_buffer[331] (data_buffer[331]), .\data_buffer[330] (data_buffer[330]), 
            .\data_buffer[329] (data_buffer[329]), .\data_buffer[328] (data_buffer[328]), 
            .\data_buffer[324] (data_buffer[324]), .\data_buffer[323] (data_buffer[323]), 
            .\data_buffer[322] (data_buffer[322]), .\data_buffer[321] (data_buffer[321]), 
            .\data_buffer[320] (data_buffer[320]), .\data_buffer[316] (data_buffer[316]), 
            .\data_buffer[315] (data_buffer[315]), .\data_buffer[314] (data_buffer[314]), 
            .\data_buffer[313] (data_buffer[313]), .\data_buffer[312] (data_buffer[312]), 
            .\data_buffer[308] (data_buffer[308]), .\data_buffer[307] (data_buffer[307]), 
            .\data_buffer[306] (data_buffer[306]), .\data_buffer[305] (data_buffer[305]), 
            .\data_buffer[304] (data_buffer[304]), .\data_buffer[300] (data_buffer[300]), 
            .\data_buffer[299] (data_buffer[299]), .\data_buffer[298] (data_buffer[298]), 
            .\data_buffer[297] (data_buffer[297]), .\data_buffer[296] (data_buffer[296]), 
            .\data_buffer[292] (data_buffer[292]), .\data_buffer[291] (data_buffer[291]), 
            .\data_buffer[290] (data_buffer[290]), .\data_buffer[289] (data_buffer[289]), 
            .\data_buffer[288] (data_buffer[288]), .\data_buffer[284] (data_buffer[284]), 
            .\data_buffer[283] (data_buffer[283]), .\data_buffer[282] (data_buffer[282]), 
            .\data_buffer[281] (data_buffer[281]), .\data_buffer[280] (data_buffer[280]), 
            .\data_buffer[276] (data_buffer[276]), .\data_buffer[275] (data_buffer[275]), 
            .\data_buffer[274] (data_buffer[274]), .\data_buffer[273] (data_buffer[273]), 
            .\data_buffer[272] (data_buffer[272]), .\data_buffer[268] (data_buffer[268]), 
            .\data_buffer[267] (data_buffer[267]), .\data_buffer[266] (data_buffer[266]), 
            .\data_buffer[265] (data_buffer[265]), .\data_buffer[264] (data_buffer[264]), 
            .\data_buffer[260] (data_buffer[260]), .\data_buffer[259] (data_buffer[259]), 
            .\data_buffer[258] (data_buffer[258]), .\data_buffer[257] (data_buffer[257]), 
            .\data_buffer[256] (data_buffer[256]), .\data_buffer[252] (data_buffer[252]), 
            .\data_buffer[251] (data_buffer[251]), .\data_buffer[250] (data_buffer[250]), 
            .\data_buffer[249] (data_buffer[249]), .\data_buffer[248] (data_buffer[248]), 
            .\data_buffer[244] (data_buffer[244]), .\data_buffer[243] (data_buffer[243]), 
            .\data_buffer[242] (data_buffer[242]), .\data_buffer[241] (data_buffer[241]), 
            .\data_buffer[240] (data_buffer[240]), .\data_buffer[236] (data_buffer[236]), 
            .\data_buffer[235] (data_buffer[235]), .\data_buffer[234] (data_buffer[234]), 
            .\data_buffer[233] (data_buffer[233]), .\data_buffer[232] (data_buffer[232]), 
            .\data_buffer[228] (data_buffer[228]), .\data_buffer[227] (data_buffer[227]), 
            .\data_buffer[226] (data_buffer[226]), .\data_buffer[225] (data_buffer[225]), 
            .\data_buffer[224] (data_buffer[224]), .\data_buffer[220] (data_buffer[220]), 
            .\data_buffer[219] (data_buffer[219]), .\data_buffer[218] (data_buffer[218]), 
            .\data_buffer[217] (data_buffer[217]), .n26793(n26793), .\data_buffer[216] (data_buffer[216]), 
            .\data_buffer[212] (data_buffer[212]), .\data_buffer[211] (data_buffer[211]), 
            .\data_buffer[210] (data_buffer[210]), .\data_buffer[209] (data_buffer[209]), 
            .\data_buffer[208] (data_buffer[208]), .\data_buffer[204] (data_buffer[204]), 
            .\data_buffer[203] (data_buffer[203]), .\data_buffer[202] (data_buffer[202]), 
            .\data_buffer[201] (data_buffer[201]), .\data_buffer[200] (data_buffer[200]), 
            .\data_buffer[196] (data_buffer[196]), .\data_buffer[195] (data_buffer[195]), 
            .\data_buffer[194] (data_buffer[194]), .\data_buffer[193] (data_buffer[193]), 
            .\data_buffer[192] (data_buffer[192]), .\data_buffer[188] (data_buffer[188]), 
            .\data_buffer[187] (data_buffer[187]), .\data_buffer[178] (data_buffer[178]), 
            .\data_buffer[170] (data_buffer[170]), .\data_buffer[179] (data_buffer[179]), 
            .\data_buffer[171] (data_buffer[171]), .\data_buffer[180] (data_buffer[180]), 
            .\data_buffer[172] (data_buffer[172]), .\data_buffer[184] (data_buffer[184]), 
            .\data_buffer[176] (data_buffer[176]), .\data_buffer[185] (data_buffer[185]), 
            .\data_buffer[177] (data_buffer[177]), .\data_buffer[186] (data_buffer[186]), 
            .\data_buffer[169] (data_buffer[169]), .\data_buffer[168] (data_buffer[168]), 
            .\data_buffer[164] (data_buffer[164]), .\data_buffer[163] (data_buffer[163]), 
            .\data_buffer[162] (data_buffer[162]), .\data_buffer[161] (data_buffer[161]), 
            .\data_buffer[160] (data_buffer[160]), .\data_buffer[156] (data_buffer[156]), 
            .\data_buffer[155] (data_buffer[155]), .\data_buffer[154] (data_buffer[154]), 
            .\data_buffer[153] (data_buffer[153]), .\data_buffer[152] (data_buffer[152]), 
            .\data_buffer[148] (data_buffer[148]), .\data_buffer[147] (data_buffer[147]), 
            .\data_buffer[146] (data_buffer[146]), .\data_buffer[145] (data_buffer[145]), 
            .\data_buffer[144] (data_buffer[144]), .\data_buffer[140] (data_buffer[140]), 
            .\data_buffer[139] (data_buffer[139]), .\data_buffer[138] (data_buffer[138]), 
            .\data_buffer[137] (data_buffer[137]), .\data_buffer[136] (data_buffer[136]), 
            .\data_buffer[132] (data_buffer[132]), .\data_buffer[131] (data_buffer[131]), 
            .\data_buffer[130] (data_buffer[130]), .\data_buffer[129] (data_buffer[129]), 
            .\data_buffer[128] (data_buffer[128]), .\data_buffer[124] (data_buffer[124]), 
            .\data_buffer[123] (data_buffer[123]), .\data_buffer[122] (data_buffer[122]), 
            .\data_buffer[121] (data_buffer[121]), .\data_buffer[120] (data_buffer[120]), 
            .\data_buffer[116] (data_buffer[116]), .\data_buffer[115] (data_buffer[115]), 
            .\data_buffer[114] (data_buffer[114]), .\data_buffer[113] (data_buffer[113]), 
            .\data_buffer[112] (data_buffer[112]), .\data_buffer[108] (data_buffer[108]), 
            .\data_buffer[107] (data_buffer[107]), .\data_buffer[106] (data_buffer[106]), 
            .\data_buffer[105] (data_buffer[105]), .\data_buffer[104] (data_buffer[104]), 
            .\data_buffer[100] (data_buffer[100]), .\data_buffer[99] (data_buffer[99]), 
            .\data_buffer[98] (data_buffer[98]), .\data_buffer[97] (data_buffer[97]), 
            .\data_buffer[96] (data_buffer[96]), .\data_buffer[92] (data_buffer[92]), 
            .\data_buffer[91] (data_buffer[91]), .\data_buffer[90] (data_buffer[90]), 
            .\data_buffer[89] (data_buffer[89]), .\data_buffer[88] (data_buffer[88]), 
            .\data_buffer[84] (data_buffer[84]), .\data_buffer[83] (data_buffer[83]), 
            .\data_buffer[82] (data_buffer[82]), .\data_buffer[81] (data_buffer[81]), 
            .\data_buffer[80] (data_buffer[80]), .\data_buffer[76] (data_buffer[76]), 
            .\data_buffer[75] (data_buffer[75]), .\data_buffer[74] (data_buffer[74]), 
            .\data_buffer[73] (data_buffer[73]), .data_length({data_length}), 
            .clk_c_enable_1399(clk_c_enable_1399), .\data_buffer[72] (data_buffer[72]), 
            .\data_buffer[68] (data_buffer[68]), .\data_buffer[67] (data_buffer[67]), 
            .\data_buffer[66] (data_buffer[66]), .\data_buffer[65] (data_buffer[65]), 
            .\data_buffer[64] (data_buffer[64]), .\data_buffer[60] (data_buffer[60]), 
            .\data_buffer[59] (data_buffer[59]), .\data_buffer[58] (data_buffer[58]), 
            .\data_buffer[57] (data_buffer[57]), .\data_buffer[56] (data_buffer[56]), 
            .\data_buffer[52] (data_buffer[52]), .\data_buffer[51] (data_buffer[51]), 
            .\data_buffer[50] (data_buffer[50]), .\data_buffer[49] (data_buffer[49]), 
            .\data_buffer[48] (data_buffer[48]), .\data_buffer[44] (data_buffer[44]), 
            .\data_buffer[43] (data_buffer[43]), .\data_buffer[42] (data_buffer[42]), 
            .\data_buffer[41] (data_buffer[41]), .\data_buffer[40] (data_buffer[40]), 
            .\data_buffer[36] (data_buffer[36]), .\data_buffer[35] (data_buffer[35]), 
            .\data_buffer[34] (data_buffer[34]), .\data_buffer[33] (data_buffer[33]), 
            .\data_buffer[32] (data_buffer[32]), .\data_buffer[28] (data_buffer[28]), 
            .\data_buffer[27] (data_buffer[27]), .\data_buffer[26] (data_buffer[26]), 
            .\data_buffer[25] (data_buffer[25]), .\data_buffer[24] (data_buffer[24]), 
            .\data_buffer[20] (data_buffer[20]), .\data_buffer[19] (data_buffer[19]), 
            .\data_buffer[18] (data_buffer[18]), .\data_buffer[17] (data_buffer[17]), 
            .\data_buffer[16] (data_buffer[16]), .\data_buffer[12] (data_buffer[12]), 
            .\data_buffer[11] (data_buffer[11]), .\data_buffer[10] (data_buffer[10]), 
            .\data_buffer[9] (data_buffer[9]), .\data_buffer[8] (data_buffer[8]), 
            .\data_buffer[4] (data_buffer[4]), .\data_buffer[3] (data_buffer[3]), 
            .\data_buffer[2] (data_buffer[2]), .\data_buffer[1] (data_buffer[1]), 
            .flag(flag), .GND_net(GND_net), .\tamp_data[0] (tamp_data[0]), 
            .\tamp_data[4] (tamp_data[4]), .\tamp_data[1] (tamp_data[1]), 
            .\tamp_data[5] (tamp_data[5]), .\tamp_data[2] (tamp_data[2]), 
            .\tamp_data[6] (tamp_data[6]), .\tamp_data[3] (tamp_data[3]), 
            .\tamp_data[7] (tamp_data[7]), .\tamp_data[9] (tamp_data[9]), 
            .\tamp_data[8] (tamp_data[8]), .n15(n15), .ready(ready), .rs232_tx_c(rs232_tx_c), 
            .rs232_rx_c(rs232_rx_c)) /* synthesis syn_module_defined=1 */ ;   // g:/fpga/mxo2/system/project/system_top.v(91[1] 101[2])
    PFUMX i22178 (.BLUT(n25806), .ALUT(n25807), .C0(cnt_adj_5212[3]), 
          .Z(n25808));
    DS18B20Z DS18B20Z_inst (.clk_1mhz(clk_1mhz), .clk_c(clk_c), .\tamp_data[0] (tamp_data[0]), 
            .clk_c_enable_931(clk_c_enable_931), .tamp_out_11__N_495(tamp_out_11__N_495), 
            .\state_back_2__N_261[2] (state_back_2__N_261[2]), .one_wire_N_501(one_wire_N_501), 
            .\state[0] (state[0]), .clk_c_enable_1439(clk_c_enable_1439), 
            .\data_out[0] (data_out[0]), .\cnt_read[2] (cnt_read[2]), .\state[1] (state[1]), 
            .\tamp_data[9] (tamp_data[9]), .\tamp_data[8] (tamp_data[8]), 
            .\tamp_data[7] (tamp_data[7]), .\tamp_data[6] (tamp_data[6]), 
            .\tamp_data[5] (tamp_data[5]), .\tamp_data[4] (tamp_data[4]), 
            .\tamp_data[2] (tamp_data[2]), .tamp_out_11__N_483(tamp_out_11__N_483), 
            .\tamp_data[1] (tamp_data[1]), .tamp_out_11__N_489(tamp_out_11__N_489), 
            .clk_c_enable_686(clk_c_enable_686), .clk_c_enable_117(clk_c_enable_117), 
            .clk_c_enable_132(clk_c_enable_132), .one_wire_out(one_wire_out), 
            .n25765(n25765), .n50(n50), .GND_net(GND_net), .n25618(n25618), 
            .n25607(n25607), .clk_c_enable_684(clk_c_enable_684), .\num_delay_19__N_369[5] (num_delay_19__N_369[5]), 
            .clk_c_enable_688(clk_c_enable_688), .\data_out[1] (data_out[1]), 
            .\data_out[2] (data_out[2]), .\tamp_out_11__N_478[3] (tamp_out_11__N_478[3]), 
            .\tamp_data[3] (tamp_data[3]), .n20945(n20945), .\cnt_init[2] (cnt_init[2]), 
            .n25689(n25689), .clk_c_enable_1433(clk_c_enable_1433), .clk_c_enable_1437(clk_c_enable_1437), 
            .n23656(n23656), .n28(n28), .n16451(n16451), .n16602(n16602), 
            .n25742(n25742), .n5709(n5709), .n37(n37), .n29(n29), .n25484(n25484), 
            .n25453(n25453), .n25857(n25857)) /* synthesis syn_module_defined=1 */ ;   // g:/fpga/mxo2/system/project/system_top.v(61[10] 67[2])
    
endmodule
//
// Verilog Description of module TSALL
// module not written out since it is a black-box. 
//

//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

//
// Verilog Description of module time_generator
//

module time_generator (time_data, clk_c, flag, n26780, en_c, key_c_1, 
            key_c_0, key_c_2, \data_out[1] , \tamp_out_11__N_478[3] , 
            \data_out[2] , tamp_out_11__N_483, \data_out[0] , tamp_out_11__N_489, 
            \data_length_reg[0] , n15, n5151, GND_net, tamp_out_11__N_495) /* synthesis syn_module_defined=1 */ ;
    output [23:0]time_data;
    input clk_c;
    output flag;
    input n26780;
    input en_c;
    input key_c_1;
    input key_c_0;
    input key_c_2;
    input \data_out[1] ;
    input \tamp_out_11__N_478[3] ;
    input \data_out[2] ;
    output tamp_out_11__N_483;
    input \data_out[0] ;
    output tamp_out_11__N_489;
    input \data_length_reg[0] ;
    input n15;
    output n5151;
    input GND_net;
    output tamp_out_11__N_495;
    
    wire clk_5hz /* synthesis is_clock=1, SET_AS_NETWORK=\time_generator_inst/clk_5hz */ ;   // g:/fpga/mxo2/system/project/time_generator.v(11[9:16])
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // g:/fpga/mxo2/system/project/system_top.v(2[15:18])
    
    wire time_out_15__N_118, n5004;
    wire [7:0]n222;
    
    wire clk_5hz_enable_11, n5006;
    wire [7:0]n280;
    wire [23:0]cnt_5hz;   // g:/fpga/mxo2/system/project/time_generator.v(12[14:21])
    
    wire clk_c_enable_682, clk_c_enable_750;
    wire [23:0]n1;
    
    wire n25724;
    wire [2:0]cnt;   // g:/fpga/mxo2/system/project/time_generator.v(23[21:24])
    
    wire cnt_2__N_88, n20922, time_out_23__N_98, n5002, n25730, n12, 
        n23131, n25725, n7, clk_c_enable_118, n22, n16, n24, n23610, 
        n20, n25726, n24024, n25664, n4, n23511, clk_5hz_enable_4;
    wire [3:0]n211;
    
    wire n24026, clk_5hz_enable_7;
    wire [3:0]n269;
    
    wire n25704, n10023, n25647, n25727, n25728, n25731, n25729;
    wire [7:0]n160;
    
    wire n24028;
    wire [3:0]n149;
    wire [2:0]n114;
    
    wire n23791, n25656, clk_5hz_enable_14, n23696, n7_adj_5193, n23805, 
        n23783, n25_adj_5194, n24044, n6, n20_adj_5195, n16_adj_5196, 
        n18_adj_5197, n20478, n20477, n20476, n20475, n20474, n20473, 
        n24_adj_5199, n23111, n20472, n23634, n20468, n20469, n20471, 
        n20467, n20470;
    
    FD1P3IX time_fen__i1 (.D(n222[0]), .SP(time_out_15__N_118), .CD(n5004), 
            .CK(clk_5hz), .Q(time_data[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=51, LSE_RLINE=58 */ ;   // g:/fpga/mxo2/system/project/time_generator.v(55[10] 64[8])
    defparam time_fen__i1.GSR = "ENABLED";
    FD1P3IX time_miao__i1 (.D(n280[0]), .SP(clk_5hz_enable_11), .CD(n5006), 
            .CK(clk_5hz), .Q(time_data[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=51, LSE_RLINE=58 */ ;   // g:/fpga/mxo2/system/project/time_generator.v(70[10] 79[8])
    defparam time_miao__i1.GSR = "ENABLED";
    FD1P3IX cnt_5hz__i0 (.D(n1[0]), .SP(clk_c_enable_682), .CD(clk_c_enable_750), 
            .CK(clk_c), .Q(cnt_5hz[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=51, LSE_RLINE=58 */ ;   // g:/fpga/mxo2/system/project/time_generator.v(16[10] 19[35])
    defparam cnt_5hz__i0.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_442 (.A(time_data[4]), .B(time_data[6]), .Z(n25724)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_442.init = 16'h8888;
    FD1S3IX cnt__i0 (.D(n20922), .CK(clk_c), .CD(cnt_2__N_88), .Q(cnt[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=51, LSE_RLINE=58 */ ;   // g:/fpga/mxo2/system/project/time_generator.v(27[10] 30[27])
    defparam cnt__i0.GSR = "ENABLED";
    FD1P3IX time_shi__i1 (.D(n25730), .SP(time_out_23__N_98), .CD(n5002), 
            .CK(clk_5hz), .Q(time_data[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=51, LSE_RLINE=58 */ ;   // g:/fpga/mxo2/system/project/time_generator.v(40[10] 49[8])
    defparam time_shi__i1.GSR = "ENABLED";
    LUT4 i5_4_lut (.A(cnt_5hz[14]), .B(cnt_5hz[23]), .C(cnt_5hz[13]), 
         .D(cnt_5hz[22]), .Z(n12)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i5_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut_3_lut_4_lut (.A(time_data[4]), .B(time_data[6]), .C(n23131), 
         .D(n25725), .Z(n7)) /* synthesis lut_function=(((C+!(D))+!B)+!A) */ ;
    defparam i2_2_lut_3_lut_4_lut.init = 16'hf7ff;
    FD1P3IX flag_100 (.D(n26780), .SP(clk_c_enable_118), .CD(flag), .CK(clk_c), 
            .Q(flag)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=51, LSE_RLINE=58 */ ;   // g:/fpga/mxo2/system/project/time_generator.v(86[10] 89[22])
    defparam flag_100.GSR = "ENABLED";
    LUT4 i11_4_lut (.A(cnt_5hz[4]), .B(n22), .C(n16), .D(cnt_5hz[1]), 
         .Z(n24)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i11_4_lut.init = 16'hfffe;
    LUT4 i7_4_lut (.A(cnt_5hz[20]), .B(cnt_5hz[11]), .C(n23610), .D(cnt_5hz[6]), 
         .Z(n20)) /* synthesis lut_function=((B+((D)+!C))+!A) */ ;
    defparam i7_4_lut.init = 16'hffdf;
    LUT4 i9_4_lut (.A(cnt_5hz[21]), .B(cnt_5hz[9]), .C(cnt_5hz[2]), .D(cnt_5hz[12]), 
         .Z(n22)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i9_4_lut.init = 16'hfffe;
    LUT4 i13389_2_lut_rep_443 (.A(time_data[0]), .B(time_data[3]), .Z(n25725)) /* synthesis lut_function=(A (B)) */ ;
    defparam i13389_2_lut_rep_443.init = 16'h8888;
    LUT4 i21309_2_lut_3_lut_4_lut (.A(time_data[0]), .B(time_data[3]), .C(time_data[4]), 
         .D(n25726), .Z(n24024)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C))+!A (C)) */ ;
    defparam i21309_2_lut_3_lut_4_lut.init = 16'hf078;
    LUT4 i3_2_lut (.A(cnt_5hz[3]), .B(cnt_5hz[0]), .Z(n16)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i3_2_lut.init = 16'heeee;
    LUT4 i20751_2_lut (.A(cnt_5hz[17]), .B(cnt_5hz[19]), .Z(n23610)) /* synthesis lut_function=(A (B)) */ ;
    defparam i20751_2_lut.init = 16'h8888;
    LUT4 en_I_0_106_4_lut (.A(en_c), .B(n25664), .C(key_c_1), .D(n4), 
         .Z(time_out_15__N_118)) /* synthesis lut_function=(!((B (C (D))+!B (C))+!A)) */ ;   // g:/fpga/mxo2/system/project/time_generator.v(55[14:99])
    defparam en_I_0_106_4_lut.init = 16'h0a8a;
    LUT4 i20675_2_lut_3_lut_4_lut (.A(time_data[0]), .B(time_data[3]), .C(time_data[5]), 
         .D(n25726), .Z(n23511)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam i20675_2_lut_3_lut_4_lut.init = 16'hfff7;
    FD1P3IX time_fen__i8 (.D(n211[3]), .SP(clk_5hz_enable_4), .CD(n5004), 
            .CK(clk_5hz), .Q(time_data[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=51, LSE_RLINE=58 */ ;   // g:/fpga/mxo2/system/project/time_generator.v(55[10] 64[8])
    defparam time_fen__i8.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_382_3_lut_4_lut (.A(time_data[0]), .B(time_data[3]), 
         .C(time_data[6]), .D(time_data[4]), .Z(n25664)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_rep_382_3_lut_4_lut.init = 16'h8000;
    FD1P3IX time_fen__i7 (.D(n211[2]), .SP(clk_5hz_enable_4), .CD(n5004), 
            .CK(clk_5hz), .Q(time_data[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=51, LSE_RLINE=58 */ ;   // g:/fpga/mxo2/system/project/time_generator.v(55[10] 64[8])
    defparam time_fen__i7.GSR = "ENABLED";
    FD1P3IX time_fen__i6 (.D(n211[1]), .SP(clk_5hz_enable_4), .CD(n5004), 
            .CK(clk_5hz), .Q(time_data[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=51, LSE_RLINE=58 */ ;   // g:/fpga/mxo2/system/project/time_generator.v(55[10] 64[8])
    defparam time_fen__i6.GSR = "ENABLED";
    FD1P3IX cnt_5hz__i23 (.D(n1[23]), .SP(clk_c_enable_682), .CD(clk_c_enable_750), 
            .CK(clk_c), .Q(cnt_5hz[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=51, LSE_RLINE=58 */ ;   // g:/fpga/mxo2/system/project/time_generator.v(16[10] 19[35])
    defparam cnt_5hz__i23.GSR = "ENABLED";
    FD1P3IX cnt_5hz__i22 (.D(n1[22]), .SP(clk_c_enable_682), .CD(clk_c_enable_750), 
            .CK(clk_c), .Q(cnt_5hz[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=51, LSE_RLINE=58 */ ;   // g:/fpga/mxo2/system/project/time_generator.v(16[10] 19[35])
    defparam cnt_5hz__i22.GSR = "ENABLED";
    FD1P3IX cnt_5hz__i21 (.D(n1[21]), .SP(clk_c_enable_682), .CD(clk_c_enable_750), 
            .CK(clk_c), .Q(cnt_5hz[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=51, LSE_RLINE=58 */ ;   // g:/fpga/mxo2/system/project/time_generator.v(16[10] 19[35])
    defparam cnt_5hz__i21.GSR = "ENABLED";
    FD1P3IX cnt_5hz__i20 (.D(n1[20]), .SP(clk_c_enable_682), .CD(clk_c_enable_750), 
            .CK(clk_c), .Q(cnt_5hz[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=51, LSE_RLINE=58 */ ;   // g:/fpga/mxo2/system/project/time_generator.v(16[10] 19[35])
    defparam cnt_5hz__i20.GSR = "ENABLED";
    FD1P3IX cnt_5hz__i19 (.D(n1[19]), .SP(clk_c_enable_682), .CD(clk_c_enable_750), 
            .CK(clk_c), .Q(cnt_5hz[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=51, LSE_RLINE=58 */ ;   // g:/fpga/mxo2/system/project/time_generator.v(16[10] 19[35])
    defparam cnt_5hz__i19.GSR = "ENABLED";
    FD1P3IX cnt_5hz__i18 (.D(n1[18]), .SP(clk_c_enable_682), .CD(clk_c_enable_750), 
            .CK(clk_c), .Q(cnt_5hz[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=51, LSE_RLINE=58 */ ;   // g:/fpga/mxo2/system/project/time_generator.v(16[10] 19[35])
    defparam cnt_5hz__i18.GSR = "ENABLED";
    FD1P3IX cnt_5hz__i17 (.D(n1[17]), .SP(clk_c_enable_682), .CD(clk_c_enable_750), 
            .CK(clk_c), .Q(cnt_5hz[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=51, LSE_RLINE=58 */ ;   // g:/fpga/mxo2/system/project/time_generator.v(16[10] 19[35])
    defparam cnt_5hz__i17.GSR = "ENABLED";
    FD1P3IX cnt_5hz__i16 (.D(n1[16]), .SP(clk_c_enable_682), .CD(clk_c_enable_750), 
            .CK(clk_c), .Q(cnt_5hz[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=51, LSE_RLINE=58 */ ;   // g:/fpga/mxo2/system/project/time_generator.v(16[10] 19[35])
    defparam cnt_5hz__i16.GSR = "ENABLED";
    FD1P3IX cnt_5hz__i15 (.D(n1[15]), .SP(clk_c_enable_682), .CD(clk_c_enable_750), 
            .CK(clk_c), .Q(cnt_5hz[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=51, LSE_RLINE=58 */ ;   // g:/fpga/mxo2/system/project/time_generator.v(16[10] 19[35])
    defparam cnt_5hz__i15.GSR = "ENABLED";
    FD1P3IX cnt_5hz__i14 (.D(n1[14]), .SP(clk_c_enable_682), .CD(clk_c_enable_750), 
            .CK(clk_c), .Q(cnt_5hz[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=51, LSE_RLINE=58 */ ;   // g:/fpga/mxo2/system/project/time_generator.v(16[10] 19[35])
    defparam cnt_5hz__i14.GSR = "ENABLED";
    FD1P3IX cnt_5hz__i13 (.D(n1[13]), .SP(clk_c_enable_682), .CD(clk_c_enable_750), 
            .CK(clk_c), .Q(cnt_5hz[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=51, LSE_RLINE=58 */ ;   // g:/fpga/mxo2/system/project/time_generator.v(16[10] 19[35])
    defparam cnt_5hz__i13.GSR = "ENABLED";
    FD1P3IX time_fen__i5 (.D(n24026), .SP(time_out_15__N_118), .CD(n5004), 
            .CK(clk_5hz), .Q(time_data[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=51, LSE_RLINE=58 */ ;   // g:/fpga/mxo2/system/project/time_generator.v(55[10] 64[8])
    defparam time_fen__i5.GSR = "ENABLED";
    FD1P3IX cnt_5hz__i12 (.D(n1[12]), .SP(clk_c_enable_682), .CD(clk_c_enable_750), 
            .CK(clk_c), .Q(cnt_5hz[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=51, LSE_RLINE=58 */ ;   // g:/fpga/mxo2/system/project/time_generator.v(16[10] 19[35])
    defparam cnt_5hz__i12.GSR = "ENABLED";
    FD1P3IX cnt_5hz__i11 (.D(n1[11]), .SP(clk_c_enable_682), .CD(clk_c_enable_750), 
            .CK(clk_c), .Q(cnt_5hz[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=51, LSE_RLINE=58 */ ;   // g:/fpga/mxo2/system/project/time_generator.v(16[10] 19[35])
    defparam cnt_5hz__i11.GSR = "ENABLED";
    FD1P3IX time_fen__i4 (.D(n222[3]), .SP(time_out_15__N_118), .CD(n5004), 
            .CK(clk_5hz), .Q(time_data[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=51, LSE_RLINE=58 */ ;   // g:/fpga/mxo2/system/project/time_generator.v(55[10] 64[8])
    defparam time_fen__i4.GSR = "ENABLED";
    FD1P3IX cnt_5hz__i10 (.D(n1[10]), .SP(clk_c_enable_682), .CD(clk_c_enable_750), 
            .CK(clk_c), .Q(cnt_5hz[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=51, LSE_RLINE=58 */ ;   // g:/fpga/mxo2/system/project/time_generator.v(16[10] 19[35])
    defparam cnt_5hz__i10.GSR = "ENABLED";
    FD1P3IX cnt_5hz__i9 (.D(n1[9]), .SP(clk_c_enable_682), .CD(clk_c_enable_750), 
            .CK(clk_c), .Q(cnt_5hz[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=51, LSE_RLINE=58 */ ;   // g:/fpga/mxo2/system/project/time_generator.v(16[10] 19[35])
    defparam cnt_5hz__i9.GSR = "ENABLED";
    FD1P3IX time_fen__i3 (.D(n222[2]), .SP(time_out_15__N_118), .CD(n5004), 
            .CK(clk_5hz), .Q(time_data[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=51, LSE_RLINE=58 */ ;   // g:/fpga/mxo2/system/project/time_generator.v(55[10] 64[8])
    defparam time_fen__i3.GSR = "ENABLED";
    FD1P3IX cnt_5hz__i8 (.D(n1[8]), .SP(clk_c_enable_682), .CD(clk_c_enable_750), 
            .CK(clk_c), .Q(cnt_5hz[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=51, LSE_RLINE=58 */ ;   // g:/fpga/mxo2/system/project/time_generator.v(16[10] 19[35])
    defparam cnt_5hz__i8.GSR = "ENABLED";
    FD1P3IX cnt_5hz__i7 (.D(n1[7]), .SP(clk_c_enable_682), .CD(clk_c_enable_750), 
            .CK(clk_c), .Q(cnt_5hz[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=51, LSE_RLINE=58 */ ;   // g:/fpga/mxo2/system/project/time_generator.v(16[10] 19[35])
    defparam cnt_5hz__i7.GSR = "ENABLED";
    FD1P3IX time_fen__i2 (.D(n222[1]), .SP(time_out_15__N_118), .CD(n5004), 
            .CK(clk_5hz), .Q(time_data[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=51, LSE_RLINE=58 */ ;   // g:/fpga/mxo2/system/project/time_generator.v(55[10] 64[8])
    defparam time_fen__i2.GSR = "ENABLED";
    FD1P3IX cnt_5hz__i6 (.D(n1[6]), .SP(clk_c_enable_682), .CD(clk_c_enable_750), 
            .CK(clk_c), .Q(cnt_5hz[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=51, LSE_RLINE=58 */ ;   // g:/fpga/mxo2/system/project/time_generator.v(16[10] 19[35])
    defparam cnt_5hz__i6.GSR = "ENABLED";
    FD1P3IX cnt_5hz__i5 (.D(n1[5]), .SP(clk_c_enable_682), .CD(clk_c_enable_750), 
            .CK(clk_c), .Q(cnt_5hz[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=51, LSE_RLINE=58 */ ;   // g:/fpga/mxo2/system/project/time_generator.v(16[10] 19[35])
    defparam cnt_5hz__i5.GSR = "ENABLED";
    FD1P3IX cnt_5hz__i4 (.D(n1[4]), .SP(clk_c_enable_682), .CD(clk_c_enable_750), 
            .CK(clk_c), .Q(cnt_5hz[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=51, LSE_RLINE=58 */ ;   // g:/fpga/mxo2/system/project/time_generator.v(16[10] 19[35])
    defparam cnt_5hz__i4.GSR = "ENABLED";
    FD1P3IX cnt_5hz__i3 (.D(n1[3]), .SP(clk_c_enable_682), .CD(clk_c_enable_750), 
            .CK(clk_c), .Q(cnt_5hz[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=51, LSE_RLINE=58 */ ;   // g:/fpga/mxo2/system/project/time_generator.v(16[10] 19[35])
    defparam cnt_5hz__i3.GSR = "ENABLED";
    FD1P3IX cnt_5hz__i2 (.D(n1[2]), .SP(clk_c_enable_682), .CD(clk_c_enable_750), 
            .CK(clk_c), .Q(cnt_5hz[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=51, LSE_RLINE=58 */ ;   // g:/fpga/mxo2/system/project/time_generator.v(16[10] 19[35])
    defparam cnt_5hz__i2.GSR = "ENABLED";
    FD1P3IX cnt_5hz__i1 (.D(n1[1]), .SP(clk_c_enable_682), .CD(clk_c_enable_750), 
            .CK(clk_c), .Q(cnt_5hz[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=51, LSE_RLINE=58 */ ;   // g:/fpga/mxo2/system/project/time_generator.v(16[10] 19[35])
    defparam cnt_5hz__i1.GSR = "ENABLED";
    FD1P3IX time_miao__i8 (.D(n269[3]), .SP(clk_5hz_enable_7), .CD(n5006), 
            .CK(clk_5hz), .Q(time_data[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=51, LSE_RLINE=58 */ ;   // g:/fpga/mxo2/system/project/time_generator.v(70[10] 79[8])
    defparam time_miao__i8.GSR = "ENABLED";
    FD1P3IX time_miao__i7 (.D(n269[2]), .SP(clk_5hz_enable_7), .CD(n5006), 
            .CK(clk_5hz), .Q(time_data[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=51, LSE_RLINE=58 */ ;   // g:/fpga/mxo2/system/project/time_generator.v(70[10] 79[8])
    defparam time_miao__i7.GSR = "ENABLED";
    FD1P3IX time_miao__i6 (.D(n269[1]), .SP(clk_5hz_enable_7), .CD(n5006), 
            .CK(clk_5hz), .Q(time_data[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=51, LSE_RLINE=58 */ ;   // g:/fpga/mxo2/system/project/time_generator.v(70[10] 79[8])
    defparam time_miao__i6.GSR = "ENABLED";
    FD1P3IX time_miao__i5 (.D(n24024), .SP(clk_5hz_enable_11), .CD(n5006), 
            .CK(clk_5hz), .Q(time_data[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=51, LSE_RLINE=58 */ ;   // g:/fpga/mxo2/system/project/time_generator.v(70[10] 79[8])
    defparam time_miao__i5.GSR = "ENABLED";
    FD1P3IX time_miao__i4 (.D(n280[3]), .SP(clk_5hz_enable_11), .CD(n5006), 
            .CK(clk_5hz), .Q(time_data[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=51, LSE_RLINE=58 */ ;   // g:/fpga/mxo2/system/project/time_generator.v(70[10] 79[8])
    defparam time_miao__i4.GSR = "ENABLED";
    FD1P3IX time_miao__i3 (.D(n280[2]), .SP(clk_5hz_enable_11), .CD(n5006), 
            .CK(clk_5hz), .Q(time_data[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=51, LSE_RLINE=58 */ ;   // g:/fpga/mxo2/system/project/time_generator.v(70[10] 79[8])
    defparam time_miao__i3.GSR = "ENABLED";
    FD1P3IX time_miao__i2 (.D(n280[1]), .SP(clk_5hz_enable_11), .CD(n5006), 
            .CK(clk_5hz), .Q(time_data[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=51, LSE_RLINE=58 */ ;   // g:/fpga/mxo2/system/project/time_generator.v(70[10] 79[8])
    defparam time_miao__i2.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_444 (.A(time_data[2]), .B(time_data[1]), .Z(n25726)) /* synthesis lut_function=(A+(B)) */ ;   // g:/fpga/mxo2/system/project/time_generator.v(88[14:28])
    defparam i1_2_lut_rep_444.init = 16'heeee;
    LUT4 en_I_0_3_lut_rep_335_4_lut (.A(cnt[2]), .B(n25704), .C(key_c_0), 
         .D(en_c), .Z(clk_5hz_enable_11)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(D))+!A (C+!(D)))) */ ;   // g:/fpga/mxo2/system/project/time_generator.v(40[116:127])
    defparam en_I_0_3_lut_rep_335_4_lut.init = 16'h2f00;
    LUT4 i2_3_lut_4_lut (.A(time_data[2]), .B(time_data[1]), .C(time_data[7]), 
         .D(time_data[5]), .Z(n10023)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // g:/fpga/mxo2/system/project/time_generator.v(88[14:28])
    defparam i2_3_lut_4_lut.init = 16'hfffe;
    LUT4 i13064_2_lut_3_lut_1_lut_1_lut (.A(time_data[0]), .Z(n280[0])) /* synthesis lut_function=(!(A)) */ ;   // g:/fpga/mxo2/system/project/time_generator.v(88[14:28])
    defparam i13064_2_lut_3_lut_1_lut_1_lut.init = 16'h5555;
    LUT4 i13227_3_lut_4_lut_4_lut_4_lut (.A(time_data[2]), .B(time_data[1]), 
         .C(time_data[3]), .D(time_data[0]), .Z(n280[1])) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A (B (D)+!B (C+!(D))))) */ ;   // g:/fpga/mxo2/system/project/time_generator.v(88[14:28])
    defparam i13227_3_lut_4_lut_4_lut_4_lut.init = 16'h23cc;
    LUT4 i1_2_lut_rep_365_3_lut_4_lut (.A(time_data[2]), .B(time_data[1]), 
         .C(time_data[3]), .D(time_data[0]), .Z(n25647)) /* synthesis lut_function=(A+(B+!(C (D)))) */ ;   // g:/fpga/mxo2/system/project/time_generator.v(88[14:28])
    defparam i1_2_lut_rep_365_3_lut_4_lut.init = 16'hefff;
    LUT4 i1_2_lut_rep_445 (.A(time_data[10]), .B(time_data[9]), .Z(n25727)) /* synthesis lut_function=(A+(B)) */ ;   // g:/fpga/mxo2/system/project/time_generator.v(40[22:41])
    defparam i1_2_lut_rep_445.init = 16'heeee;
    LUT4 i21582_2_lut_2_lut_3_lut_4_lut (.A(time_data[10]), .B(time_data[9]), 
         .C(time_out_15__N_118), .D(n25728), .Z(clk_5hz_enable_4)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // g:/fpga/mxo2/system/project/time_generator.v(40[22:41])
    defparam i21582_2_lut_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i21311_2_lut_3_lut_4_lut (.A(time_data[10]), .B(time_data[9]), 
         .C(time_data[12]), .D(n25728), .Z(n24026)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !(C (D)+!C !(D)))) */ ;   // g:/fpga/mxo2/system/project/time_generator.v(40[22:41])
    defparam i21311_2_lut_3_lut_4_lut.init = 16'he1f0;
    LUT4 i13358_2_lut_rep_446 (.A(time_data[8]), .B(time_data[11]), .Z(n25728)) /* synthesis lut_function=(A (B)) */ ;
    defparam i13358_2_lut_rep_446.init = 16'h8888;
    LUT4 i13289_4_lut (.A(time_data[19]), .B(n25731), .C(time_data[18]), 
         .D(n25729), .Z(n160[3])) /* synthesis lut_function=(!(A ((C (D))+!B)+!A !(B (C (D))))) */ ;   // g:/fpga/mxo2/system/project/time_generator.v(48[13:51])
    defparam i13289_4_lut.init = 16'h4888;
    LUT4 i21313_2_lut (.A(time_data[20]), .B(n25731), .Z(n24028)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // g:/fpga/mxo2/system/project/time_generator.v(48[13:51])
    defparam i21313_2_lut.init = 16'h9999;
    LUT4 i2433_2_lut (.A(time_data[21]), .B(time_data[20]), .Z(n149[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // g:/fpga/mxo2/system/project/time_generator.v(44[30:50])
    defparam i2433_2_lut.init = 16'h6666;
    LUT4 i13061_2_lut_3_lut_4_lut_1_lut (.A(time_data[8]), .Z(n222[0])) /* synthesis lut_function=(!(A)) */ ;
    defparam i13061_2_lut_3_lut_4_lut_1_lut.init = 16'h5555;
    LUT4 i13233_3_lut_4_lut_4_lut_4_lut (.A(time_data[8]), .B(time_data[11]), 
         .C(time_data[9]), .D(time_data[10]), .Z(n222[1])) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C))+!A !(C))) */ ;
    defparam i13233_3_lut_4_lut_4_lut_4_lut.init = 16'h5a52;
    FD1P3IX cnt__i1 (.D(n114[1]), .SP(clk_c_enable_750), .CD(cnt_2__N_88), 
            .CK(clk_c), .Q(cnt[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=51, LSE_RLINE=58 */ ;   // g:/fpga/mxo2/system/project/time_generator.v(27[10] 30[27])
    defparam cnt__i1.GSR = "ENABLED";
    FD1P3IX cnt__i2 (.D(n114[2]), .SP(clk_c_enable_750), .CD(cnt_2__N_88), 
            .CK(clk_c), .Q(cnt[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=51, LSE_RLINE=58 */ ;   // g:/fpga/mxo2/system/project/time_generator.v(27[10] 30[27])
    defparam cnt__i2.GSR = "ENABLED";
    LUT4 i3_4_lut (.A(time_data[14]), .B(time_data[12]), .C(time_out_15__N_118), 
         .D(n23791), .Z(n5004)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i3_4_lut.init = 16'h0080;
    LUT4 i21569_2_lut_2_lut_4_lut (.A(en_c), .B(n25656), .C(key_c_0), 
         .D(n25647), .Z(clk_5hz_enable_7)) /* synthesis lut_function=(!((B (C+(D))+!B (D))+!A)) */ ;   // g:/fpga/mxo2/system/project/time_generator.v(70[15:49])
    defparam i21569_2_lut_2_lut_4_lut.init = 16'h002a;
    LUT4 i2464_2_lut_rep_447 (.A(time_data[17]), .B(time_data[16]), .Z(n25729)) /* synthesis lut_function=(A (B)) */ ;   // g:/fpga/mxo2/system/project/time_generator.v(48[30:50])
    defparam i2464_2_lut_rep_447.init = 16'h8888;
    LUT4 i2460_1_lut_rep_448 (.A(time_data[16]), .Z(n25730)) /* synthesis lut_function=(!(A)) */ ;   // g:/fpga/mxo2/system/project/time_generator.v(48[30:50])
    defparam i2460_1_lut_rep_448.init = 16'h5555;
    LUT4 i3_4_lut_rep_449 (.A(time_data[16]), .B(time_data[19]), .C(time_data[17]), 
         .D(time_data[18]), .Z(n25731)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;   // g:/fpga/mxo2/system/project/time_generator.v(48[30:50])
    defparam i3_4_lut_rep_449.init = 16'hfff7;
    LUT4 i13292_3_lut_4_lut (.A(time_data[16]), .B(time_data[19]), .C(time_data[17]), 
         .D(time_data[18]), .Z(n160[1])) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C))+!A !(C))) */ ;   // g:/fpga/mxo2/system/project/time_generator.v(48[30:50])
    defparam i13292_3_lut_4_lut.init = 16'h5a52;
    LUT4 i13291_3_lut_4_lut_3_lut (.A(time_data[16]), .B(time_data[17]), 
         .C(time_data[18]), .Z(n160[2])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // g:/fpga/mxo2/system/project/time_generator.v(48[30:50])
    defparam i13291_3_lut_4_lut_3_lut.init = 16'h7878;
    FD1P3IX time_shi__i2 (.D(n160[1]), .SP(time_out_23__N_98), .CD(n5002), 
            .CK(clk_5hz), .Q(time_data[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=51, LSE_RLINE=58 */ ;   // g:/fpga/mxo2/system/project/time_generator.v(40[10] 49[8])
    defparam time_shi__i2.GSR = "ENABLED";
    FD1P3IX time_shi__i3 (.D(n160[2]), .SP(time_out_23__N_98), .CD(n5002), 
            .CK(clk_5hz), .Q(time_data[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=51, LSE_RLINE=58 */ ;   // g:/fpga/mxo2/system/project/time_generator.v(40[10] 49[8])
    defparam time_shi__i3.GSR = "ENABLED";
    FD1P3IX time_shi__i4 (.D(n160[3]), .SP(time_out_23__N_98), .CD(n5002), 
            .CK(clk_5hz), .Q(time_data[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=51, LSE_RLINE=58 */ ;   // g:/fpga/mxo2/system/project/time_generator.v(40[10] 49[8])
    defparam time_shi__i4.GSR = "ENABLED";
    FD1P3IX time_shi__i5 (.D(n24028), .SP(time_out_23__N_98), .CD(n5002), 
            .CK(clk_5hz), .Q(time_data[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=51, LSE_RLINE=58 */ ;   // g:/fpga/mxo2/system/project/time_generator.v(40[10] 49[8])
    defparam time_shi__i5.GSR = "ENABLED";
    FD1P3IX time_shi__i6 (.D(n149[1]), .SP(clk_5hz_enable_14), .CD(n5002), 
            .CK(clk_5hz), .Q(time_data[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=51, LSE_RLINE=58 */ ;   // g:/fpga/mxo2/system/project/time_generator.v(40[10] 49[8])
    defparam time_shi__i6.GSR = "ENABLED";
    FD1P3IX time_shi__i7 (.D(n149[2]), .SP(clk_5hz_enable_14), .CD(n5002), 
            .CK(clk_5hz), .Q(time_data[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=51, LSE_RLINE=58 */ ;   // g:/fpga/mxo2/system/project/time_generator.v(40[10] 49[8])
    defparam time_shi__i7.GSR = "ENABLED";
    FD1P3IX time_shi__i8 (.D(n149[3]), .SP(clk_5hz_enable_14), .CD(n5002), 
            .CK(clk_5hz), .Q(time_data[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=51, LSE_RLINE=58 */ ;   // g:/fpga/mxo2/system/project/time_generator.v(40[10] 49[8])
    defparam time_shi__i8.GSR = "ENABLED";
    LUT4 en_I_0_104_4_lut (.A(en_c), .B(n7), .C(key_c_2), .D(n23696), 
         .Z(time_out_23__N_98)) /* synthesis lut_function=(!((B (C)+!B !((D)+!C))+!A)) */ ;   // g:/fpga/mxo2/system/project/time_generator.v(40[14:144])
    defparam en_I_0_104_4_lut.init = 16'h2a0a;
    LUT4 i20832_4_lut (.A(time_data[12]), .B(cnt[2]), .C(time_data[14]), 
         .D(n25728), .Z(n23696)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i20832_4_lut.init = 16'h8000;
    LUT4 i5_4_lut_adj_280 (.A(time_data[21]), .B(n7_adj_5193), .C(n23805), 
         .D(n25729), .Z(n5002)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i5_4_lut_adj_280.init = 16'h0800;
    LUT4 i1_2_lut (.A(time_data[19]), .B(time_out_23__N_98), .Z(n7_adj_5193)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut.init = 16'h4444;
    LUT4 i20929_4_lut (.A(time_data[20]), .B(time_data[18]), .C(time_data[22]), 
         .D(time_data[23]), .Z(n23805)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20929_4_lut.init = 16'hfffe;
    LUT4 i21464_2_lut_4_lut_4_lut (.A(n25656), .B(n23783), .C(n25_adj_5194), 
         .D(n24044), .Z(cnt_2__N_88)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // g:/fpga/mxo2/system/project/time_generator.v(40[116:127])
    defparam i21464_2_lut_4_lut_4_lut.init = 16'h0400;
    LUT4 i4_4_lut (.A(n25727), .B(n10023), .C(time_data[15]), .D(n6), 
         .Z(n23131)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // g:/fpga/mxo2/system/project/time_generator.v(40[116:127])
    defparam i4_4_lut.init = 16'hfffe;
    LUT4 i16608_3_lut (.A(\data_out[1] ), .B(\tamp_out_11__N_478[3] ), .C(\data_out[2] ), 
         .Z(tamp_out_11__N_483)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A ((C)+!B))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(7[22:30])
    defparam i16608_3_lut.init = 16'h2c2c;
    LUT4 i16602_4_lut (.A(\data_out[2] ), .B(\data_out[0] ), .C(\tamp_out_11__N_478[3] ), 
         .D(\data_out[1] ), .Z(tamp_out_11__N_489)) /* synthesis lut_function=(!(A (C+(D))+!A !(B (C+(D))+!B (C (D))))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(7[22:30])
    defparam i16602_4_lut.init = 16'h544a;
    LUT4 i2_4_lut (.A(n25724), .B(clk_5hz_enable_11), .C(time_data[7]), 
         .D(n23511), .Z(n5006)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i2_4_lut.init = 16'h0008;
    LUT4 i2396_3_lut_4_lut (.A(time_data[5]), .B(time_data[4]), .C(time_data[6]), 
         .D(time_data[7]), .Z(n269[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // g:/fpga/mxo2/system/project/time_generator.v(74[31:52])
    defparam i2396_3_lut_4_lut.init = 16'h7f80;
    LUT4 i2389_2_lut_3_lut (.A(time_data[5]), .B(time_data[4]), .C(time_data[6]), 
         .Z(n269[2])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // g:/fpga/mxo2/system/project/time_generator.v(74[31:52])
    defparam i2389_2_lut_3_lut.init = 16'h7878;
    LUT4 i2782_3_lut_4_lut (.A(time_data[13]), .B(time_data[12]), .C(time_data[14]), 
         .D(time_data[15]), .Z(n211[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // g:/fpga/mxo2/system/project/time_generator.v(59[30:50])
    defparam i2782_3_lut_4_lut.init = 16'h7f80;
    LUT4 i2775_2_lut_3_lut (.A(time_data[13]), .B(time_data[12]), .C(time_data[14]), 
         .Z(n211[2])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // g:/fpga/mxo2/system/project/time_generator.v(59[30:50])
    defparam i2775_2_lut_3_lut.init = 16'h7878;
    LUT4 i2411_2_lut (.A(cnt[1]), .B(cnt[0]), .Z(n114[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // g:/fpga/mxo2/system/project/time_generator.v(30[16:26])
    defparam i2411_2_lut.init = 16'h6666;
    LUT4 i2418_3_lut (.A(cnt[2]), .B(cnt[1]), .C(cnt[0]), .Z(n114[2])) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;   // g:/fpga/mxo2/system/project/time_generator.v(30[16:26])
    defparam i2418_3_lut.init = 16'h6a6a;
    LUT4 i21480_4_lut (.A(time_data[11]), .B(n20_adj_5195), .C(n16_adj_5196), 
         .D(time_data[6]), .Z(clk_c_enable_118)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // g:/fpga/mxo2/system/project/time_generator.v(88[14:28])
    defparam i21480_4_lut.init = 16'h0001;
    LUT4 i9_4_lut_adj_281 (.A(clk_c_enable_750), .B(n18_adj_5197), .C(time_data[14]), 
         .D(time_data[4]), .Z(n20_adj_5195)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // g:/fpga/mxo2/system/project/time_generator.v(40[116:127])
    defparam i9_4_lut_adj_281.init = 16'hfffd;
    LUT4 i5_2_lut (.A(time_data[3]), .B(n23131), .Z(n16_adj_5196)) /* synthesis lut_function=(A+(B)) */ ;   // g:/fpga/mxo2/system/project/time_generator.v(40[116:127])
    defparam i5_2_lut.init = 16'heeee;
    LUT4 i7_4_lut_adj_282 (.A(time_data[12]), .B(cnt[2]), .C(time_data[0]), 
         .D(time_data[8]), .Z(n18_adj_5197)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // g:/fpga/mxo2/system/project/time_generator.v(40[116:127])
    defparam i7_4_lut_adj_282.init = 16'hfffe;
    LUT4 i21606_2_lut_2_lut (.A(n25731), .B(time_out_23__N_98), .Z(clk_5hz_enable_14)) /* synthesis lut_function=(!(A+!(B))) */ ;   // g:/fpga/mxo2/system/project/time_generator.v(40[10] 49[8])
    defparam i21606_2_lut_2_lut.init = 16'h4444;
    LUT4 i1_2_lut_rep_422 (.A(cnt[1]), .B(cnt[0]), .Z(n25704)) /* synthesis lut_function=(A+(B)) */ ;   // g:/fpga/mxo2/system/project/time_generator.v(40[116:127])
    defparam i1_2_lut_rep_422.init = 16'heeee;
    LUT4 i1_2_lut_3_lut (.A(cnt[1]), .B(cnt[0]), .C(time_data[13]), .Z(n6)) /* synthesis lut_function=(A+(B+(C))) */ ;   // g:/fpga/mxo2/system/project/time_generator.v(40[116:127])
    defparam i1_2_lut_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_3_lut_4_lut (.A(cnt[1]), .B(cnt[0]), .C(n10023), .D(cnt[2]), 
         .Z(n4)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // g:/fpga/mxo2/system/project/time_generator.v(40[116:127])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfeff;
    LUT4 i1_2_lut_rep_374_3_lut (.A(cnt[1]), .B(cnt[0]), .C(cnt[2]), .Z(n25656)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // g:/fpga/mxo2/system/project/time_generator.v(40[116:127])
    defparam i1_2_lut_rep_374_3_lut.init = 16'hefef;
    LUT4 i1_4_lut (.A(flag), .B(en_c), .C(\data_length_reg[0] ), .D(n15), 
         .Z(n5151)) /* synthesis lut_function=(!(A+!(B+!((D)+!C)))) */ ;   // g:/fpga/mxo2/system/project/time_generator.v(86[10] 89[22])
    defparam i1_4_lut.init = 16'h4454;
    CCU2D add_6_25 (.A0(cnt_5hz[23]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n20478), 
          .S0(n1[23]));   // g:/fpga/mxo2/system/project/time_generator.v(19[20:34])
    defparam add_6_25.INIT0 = 16'h5aaa;
    defparam add_6_25.INIT1 = 16'h0000;
    defparam add_6_25.INJECT1_0 = "NO";
    defparam add_6_25.INJECT1_1 = "NO";
    LUT4 i2768_2_lut (.A(time_data[13]), .B(time_data[12]), .Z(n211[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // g:/fpga/mxo2/system/project/time_generator.v(59[30:50])
    defparam i2768_2_lut.init = 16'h6666;
    CCU2D add_6_23 (.A0(cnt_5hz[21]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt_5hz[22]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n20477), .COUT(n20478), .S0(n1[21]), .S1(n1[22]));   // g:/fpga/mxo2/system/project/time_generator.v(19[20:34])
    defparam add_6_23.INIT0 = 16'h5aaa;
    defparam add_6_23.INIT1 = 16'h5aaa;
    defparam add_6_23.INJECT1_0 = "NO";
    defparam add_6_23.INJECT1_1 = "NO";
    CCU2D add_6_21 (.A0(cnt_5hz[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt_5hz[20]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n20476), .COUT(n20477), .S0(n1[19]), .S1(n1[20]));   // g:/fpga/mxo2/system/project/time_generator.v(19[20:34])
    defparam add_6_21.INIT0 = 16'h5aaa;
    defparam add_6_21.INIT1 = 16'h5aaa;
    defparam add_6_21.INJECT1_0 = "NO";
    defparam add_6_21.INJECT1_1 = "NO";
    CCU2D add_6_19 (.A0(cnt_5hz[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt_5hz[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n20475), .COUT(n20476), .S0(n1[17]), .S1(n1[18]));   // g:/fpga/mxo2/system/project/time_generator.v(19[20:34])
    defparam add_6_19.INIT0 = 16'h5aaa;
    defparam add_6_19.INIT1 = 16'h5aaa;
    defparam add_6_19.INJECT1_0 = "NO";
    defparam add_6_19.INJECT1_1 = "NO";
    LUT4 tamp_out_11__N_478_3__bdd_4_lut (.A(\tamp_out_11__N_478[3] ), .B(\data_out[2] ), 
         .C(\data_out[1] ), .D(\data_out[0] ), .Z(tamp_out_11__N_495)) /* synthesis lut_function=(A (B (C)+!B (C (D)+!C !(D)))+!A !(B (C)+!B (C (D)+!C !(D)))) */ ;
    defparam tamp_out_11__N_478_3__bdd_4_lut.init = 16'ha596;
    CCU2D add_6_17 (.A0(cnt_5hz[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt_5hz[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n20474), .COUT(n20475), .S0(n1[15]), .S1(n1[16]));   // g:/fpga/mxo2/system/project/time_generator.v(19[20:34])
    defparam add_6_17.INIT0 = 16'h5aaa;
    defparam add_6_17.INIT1 = 16'h5aaa;
    defparam add_6_17.INJECT1_0 = "NO";
    defparam add_6_17.INJECT1_1 = "NO";
    CCU2D add_6_15 (.A0(cnt_5hz[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt_5hz[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n20473), .COUT(n20474), .S0(n1[13]), .S1(n1[14]));   // g:/fpga/mxo2/system/project/time_generator.v(19[20:34])
    defparam add_6_15.INIT0 = 16'h5aaa;
    defparam add_6_15.INIT1 = 16'h5aaa;
    defparam add_6_15.INJECT1_0 = "NO";
    defparam add_6_15.INJECT1_1 = "NO";
    LUT4 i2382_2_lut (.A(time_data[5]), .B(time_data[4]), .Z(n269[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // g:/fpga/mxo2/system/project/time_generator.v(74[31:52])
    defparam i2382_2_lut.init = 16'h6666;
    LUT4 i13225_4_lut_4_lut (.A(time_data[3]), .B(time_data[2]), .C(time_data[1]), 
         .D(time_data[0]), .Z(n280[3])) /* synthesis lut_function=(!(A (B (C (D))+!B !(C+!(D)))+!A !(B (C (D))))) */ ;   // g:/fpga/mxo2/system/project/time_generator.v(78[13:53])
    defparam i13225_4_lut_4_lut.init = 16'h68aa;
    LUT4 i13231_4_lut_4_lut (.A(time_data[11]), .B(time_data[8]), .C(time_data[9]), 
         .D(time_data[10]), .Z(n222[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D)))+!A !(B (C (D))))) */ ;   // g:/fpga/mxo2/system/project/time_generator.v(63[13:51])
    defparam i13231_4_lut_4_lut.init = 16'h6aa2;
    LUT4 i21331_3_lut_rep_301 (.A(n24044), .B(n25_adj_5194), .C(n23783), 
         .Z(clk_c_enable_750)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // g:/fpga/mxo2/system/project/time_generator.v(88[58:80])
    defparam i21331_3_lut_rep_301.init = 16'h2020;
    LUT4 i20915_3_lut_4_lut (.A(n25727), .B(n25728), .C(time_data[13]), 
         .D(time_data[15]), .Z(n23791)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // g:/fpga/mxo2/system/project/time_generator.v(40[22:41])
    defparam i20915_3_lut_4_lut.init = 16'hfffb;
    LUT4 i1_2_lut_4_lut (.A(n24044), .B(n25_adj_5194), .C(n23783), .D(cnt[0]), 
         .Z(n20922)) /* synthesis lut_function=(A (B (D)+!B !(C (D)+!C !(D)))+!A (D)) */ ;   // g:/fpga/mxo2/system/project/time_generator.v(88[58:80])
    defparam i1_2_lut_4_lut.init = 16'hdf20;
    LUT4 i2217_2_lut_4_lut (.A(n24044), .B(n25_adj_5194), .C(n23783), 
         .D(en_c), .Z(clk_c_enable_682)) /* synthesis lut_function=(A (B (D)+!B (C+(D)))+!A (D)) */ ;   // g:/fpga/mxo2/system/project/time_generator.v(88[58:80])
    defparam i2217_2_lut_4_lut.init = 16'hff20;
    LUT4 i13232_3_lut_4_lut_4_lut_4_lut (.A(time_data[10]), .B(time_data[9]), 
         .C(time_data[8]), .Z(n222[2])) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;   // g:/fpga/mxo2/system/project/time_generator.v(40[22:41])
    defparam i13232_3_lut_4_lut_4_lut_4_lut.init = 16'h6a6a;
    LUT4 i13226_3_lut_4_lut_4_lut_4_lut (.A(time_data[2]), .B(time_data[1]), 
         .C(time_data[0]), .Z(n280[2])) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;   // g:/fpga/mxo2/system/project/time_generator.v(88[14:28])
    defparam i13226_3_lut_4_lut_4_lut_4_lut.init = 16'h6a6a;
    LUT4 i21329_4_lut (.A(cnt_5hz[1]), .B(n24_adj_5199), .C(cnt_5hz[12]), 
         .D(cnt_5hz[21]), .Z(n24044)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // g:/fpga/mxo2/system/project/time_generator.v(88[58:80])
    defparam i21329_4_lut.init = 16'h2000;
    LUT4 i10_4_lut (.A(cnt_5hz[17]), .B(n23111), .C(cnt_5hz[20]), .D(cnt_5hz[6]), 
         .Z(n25_adj_5194)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;
    defparam i10_4_lut.init = 16'hfeff;
    CCU2D add_6_13 (.A0(cnt_5hz[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt_5hz[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n20472), .COUT(n20473), .S0(n1[11]), .S1(n1[12]));   // g:/fpga/mxo2/system/project/time_generator.v(19[20:34])
    defparam add_6_13.INIT0 = 16'h5aaa;
    defparam add_6_13.INIT1 = 16'h5aaa;
    defparam add_6_13.INJECT1_0 = "NO";
    defparam add_6_13.INJECT1_1 = "NO";
    LUT4 i20907_4_lut (.A(cnt_5hz[11]), .B(cnt_5hz[2]), .C(cnt_5hz[3]), 
         .D(cnt_5hz[5]), .Z(n23783)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i20907_4_lut.init = 16'h8000;
    LUT4 i9_4_lut_adj_283 (.A(cnt_5hz[19]), .B(cnt_5hz[0]), .C(cnt_5hz[4]), 
         .D(cnt_5hz[9]), .Z(n24_adj_5199)) /* synthesis lut_function=(A+!(B (C (D)))) */ ;
    defparam i9_4_lut_adj_283.init = 16'hbfff;
    LUT4 i6_4_lut (.A(n23634), .B(n12), .C(cnt_5hz[8]), .D(cnt_5hz[16]), 
         .Z(n23111)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i6_4_lut.init = 16'hfffd;
    CCU2D add_6_5 (.A0(cnt_5hz[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt_5hz[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n20468), .COUT(n20469), .S0(n1[3]), .S1(n1[4]));   // g:/fpga/mxo2/system/project/time_generator.v(19[20:34])
    defparam add_6_5.INIT0 = 16'h5aaa;
    defparam add_6_5.INIT1 = 16'h5aaa;
    defparam add_6_5.INJECT1_0 = "NO";
    defparam add_6_5.INJECT1_1 = "NO";
    LUT4 i21483_4_lut (.A(cnt_5hz[5]), .B(n24), .C(n20), .D(n23111), 
         .Z(clk_5hz)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // g:/fpga/mxo2/system/project/time_generator.v(21[18:42])
    defparam i21483_4_lut.init = 16'h0001;
    LUT4 i2440_2_lut_3_lut (.A(time_data[21]), .B(time_data[20]), .C(time_data[22]), 
         .Z(n149[2])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // g:/fpga/mxo2/system/project/time_generator.v(44[30:50])
    defparam i2440_2_lut_3_lut.init = 16'h7878;
    CCU2D add_6_11 (.A0(cnt_5hz[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt_5hz[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n20471), .COUT(n20472), .S0(n1[9]), .S1(n1[10]));   // g:/fpga/mxo2/system/project/time_generator.v(19[20:34])
    defparam add_6_11.INIT0 = 16'h5aaa;
    defparam add_6_11.INIT1 = 16'h5aaa;
    defparam add_6_11.INJECT1_0 = "NO";
    defparam add_6_11.INJECT1_1 = "NO";
    LUT4 i2447_3_lut_4_lut (.A(time_data[21]), .B(time_data[20]), .C(time_data[22]), 
         .D(time_data[23]), .Z(n149[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // g:/fpga/mxo2/system/project/time_generator.v(44[30:50])
    defparam i2447_3_lut_4_lut.init = 16'h7f80;
    CCU2D add_6_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt_5hz[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n20467), .S1(n1[0]));   // g:/fpga/mxo2/system/project/time_generator.v(19[20:34])
    defparam add_6_1.INIT0 = 16'hF000;
    defparam add_6_1.INIT1 = 16'h5555;
    defparam add_6_1.INJECT1_0 = "NO";
    defparam add_6_1.INJECT1_1 = "NO";
    CCU2D add_6_3 (.A0(cnt_5hz[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt_5hz[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n20467), .COUT(n20468), .S0(n1[1]), .S1(n1[2]));   // g:/fpga/mxo2/system/project/time_generator.v(19[20:34])
    defparam add_6_3.INIT0 = 16'h5aaa;
    defparam add_6_3.INIT1 = 16'h5aaa;
    defparam add_6_3.INJECT1_0 = "NO";
    defparam add_6_3.INJECT1_1 = "NO";
    CCU2D add_6_9 (.A0(cnt_5hz[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt_5hz[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n20470), .COUT(n20471), .S0(n1[7]), .S1(n1[8]));   // g:/fpga/mxo2/system/project/time_generator.v(19[20:34])
    defparam add_6_9.INIT0 = 16'h5aaa;
    defparam add_6_9.INIT1 = 16'h5aaa;
    defparam add_6_9.INJECT1_0 = "NO";
    defparam add_6_9.INJECT1_1 = "NO";
    LUT4 i20773_4_lut (.A(cnt_5hz[10]), .B(cnt_5hz[15]), .C(cnt_5hz[18]), 
         .D(cnt_5hz[7]), .Z(n23634)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i20773_4_lut.init = 16'h8000;
    CCU2D add_6_7 (.A0(cnt_5hz[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt_5hz[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n20469), .COUT(n20470), .S0(n1[5]), .S1(n1[6]));   // g:/fpga/mxo2/system/project/time_generator.v(19[20:34])
    defparam add_6_7.INIT0 = 16'h5aaa;
    defparam add_6_7.INIT1 = 16'h5aaa;
    defparam add_6_7.INJECT1_0 = "NO";
    defparam add_6_7.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module OLED12832
//

module OLED12832 (clk_c, oled_csn_c, n25808, n1358, n1359, n1138, 
            n1278, n998, n579, n719, n439, n578, n718, n438, 
            n1357, n1356, n23966, n23967, cnt, n1141, n1281, n1140, 
            n1280, time_data, \tamp_data[1] , n865, n582, n722, 
            n581, n721, n1139, n1279, n999, n583, n723, n580, 
            n720, n1142, n1282, n1424, n1144, n1284, n1143, n1283, 
            n584, n724, n1355, n25751, n1354, n23974, n23971, 
            n22685, GND_net, n25774, \tamp_data[3] , n25685, n863, 
            n1423, n1425, \tamp_data[0] , \tamp_data[8] , \tamp_data[4] , 
            \tamp_data[6] , n864, oled_dat_c, n25826, oled_clk_c, 
            oled_dcn_c, \tamp_data[7] , \tamp_data[9] , \tamp_data[5] , 
            oled_rst_c, \tamp_data[2] , n1145, n585, n725, n1285) /* synthesis syn_module_defined=1 */ ;
    input clk_c;
    output oled_csn_c;
    input n25808;
    output n1358;
    output n1359;
    input n1138;
    input n1278;
    input n998;
    input n579;
    input n719;
    input n439;
    input n578;
    input n718;
    input n438;
    output n1357;
    output n1356;
    input n23966;
    input n23967;
    output [15:0]cnt;
    input n1141;
    input n1281;
    input n1140;
    input n1280;
    input [23:0]time_data;
    input \tamp_data[1] ;
    input n865;
    input n582;
    input n722;
    input n581;
    input n721;
    input n1139;
    input n1279;
    input n999;
    input n583;
    input n723;
    input n580;
    input n720;
    input n1142;
    input n1282;
    input n1424;
    input n1144;
    input n1284;
    input n1143;
    input n1283;
    input n584;
    input n724;
    output n1355;
    input n25751;
    output n1354;
    input n23974;
    input n23971;
    input n22685;
    input GND_net;
    input n25774;
    input \tamp_data[3] ;
    output n25685;
    input n863;
    input n1423;
    input n1425;
    input \tamp_data[0] ;
    input \tamp_data[8] ;
    input \tamp_data[4] ;
    input \tamp_data[6] ;
    input n864;
    output oled_dat_c;
    input n25826;
    output oled_clk_c;
    output oled_dcn_c;
    input \tamp_data[7] ;
    input \tamp_data[9] ;
    input \tamp_data[5] ;
    output oled_rst_c;
    input \tamp_data[2] ;
    input n1145;
    input n585;
    input n725;
    input n1285;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // g:/fpga/mxo2/system/project/system_top.v(2[15:18])
    wire [5:0]state;   // g:/fpga/mxo2/system/project/oled12832.v(29[13:18])
    
    wire n8, n25637;
    wire [7:0]char_reg;   // g:/fpga/mxo2/system/project/oled12832.v(26[25:33])
    wire [4:0]cnt_write;   // g:/fpga/mxo2/system/project/oled12832.v(27[43:52])
    
    wire n23877, n25635, n25630, n23422, n25601, n17, n32, n37;
    wire [4:0]cnt_main;   // g:/fpga/mxo2/system/project/oled12832.v(27[13:21])
    
    wire n43;
    wire [15:0]cnt_delay;   // g:/fpga/mxo2/system/project/oled12832.v(28[25:34])
    
    wire clk_c_enable_1452, n12055;
    wire [15:0]n2559;
    wire [4:0]cnt_init;   // g:/fpga/mxo2/system/project/oled12832.v(27[23:31])
    
    wire clk_c_enable_1359;
    wire [4:0]n3871;
    wire [7:0]y_ph;   // g:/fpga/mxo2/system/project/oled12832.v(24[16:20])
    
    wire clk_c_enable_690;
    wire [1:0]n5820;
    
    wire clk_c_enable_702;
    wire [7:0]n3492;
    wire [15:0]num1_delay;   // g:/fpga/mxo2/system/project/oled12832.v(28[13:23])
    wire [15:0]num1_delay_15__N_605;
    wire [5:0]state_back;   // g:/fpga/mxo2/system/project/oled12832.v(29[20:30])
    wire [5:0]state_back_5__N_659;
    
    wire clk_c_enable_10;
    wire [0:0]n3153;
    wire [4:0]n1;
    wire [7:0]x_ph;   // g:/fpga/mxo2/system/project/oled12832.v(23[13:17])
    wire [7:0]x_ph_7__N_519;
    
    wire n9, n25587, clk_c_enable_1352, n16632, clk_c_enable_114, 
        n25374, n25371, n25574, n23953, n16666, n25373, n25372, 
        n36, n25610, n5, n25561, n25369;
    wire [4:0]cnt_scan;   // g:/fpga/mxo2/system/project/oled12832.v(27[33:41])
    
    wire n16, n20791, n3599, n23876, n23875, n29, n16393, n9173, 
        clk_c_enable_1431;
    wire [7:0]num2;   // g:/fpga/mxo2/system/project/oled12832.v(26[19:23])
    
    wire n12049;
    wire [7:0]num2_7__N_748;
    wire [7:0]num1;   // g:/fpga/mxo2/system/project/oled12832.v(26[13:17])
    
    wire clk_c_enable_1432, n14556;
    wire [7:0]num1_7__N_732;
    wire [7:0]y_pl;   // g:/fpga/mxo2/system/project/oled12832.v(24[22:26])
    
    wire n16636, clk_c_enable_1446, n12042;
    wire [4:0]cnt_scan_4__N_682;
    
    wire n12039;
    wire [4:0]n2;
    
    wire n25558, n25038, n25040, n23134, n25557, n9304, n322, 
        n25469, n25676, n15, n25696, n25823, n23311, n21, n23, 
        n9872, n20744, n59, n41, n25682, n25638, n34, n102, 
        n80, n99, n23763, n25311, n25651, oled_dcn_N_888, n25755, 
        n23579, n23581, n23583, n25753, n25120, n25495, n8855, 
        n12, n11, n9_adj_5037, n8_adj_5038, n25800, n25801, n9_adj_5039, 
        n8_adj_5040, n23415, n31, n25325, n25323, n25326, n25553, 
        n25686, n25519, n15_adj_5041, n25650, n23253, n12_adj_5042, 
        n25599, n25566, n92, n10074, n25315, n25314, n25316, n12_adj_5043, 
        n25621, n22121, n17_adj_5044, clk_c_enable_1374, n42, n46, 
        n12_adj_5045, n25312, n25313, n25537, n23694, n25586, n23281, 
        n23347, n25632, n23348, n25538, n9_adj_5046;
    wire [7:0]char;   // g:/fpga/mxo2/system/project/oled12832.v(25[13:17])
    
    wire n25785, n9_adj_5047, n68, n69, n7, n4, n5_adj_5048, n6, 
        n23879, n23880, n23881, n12_adj_5049, n11_adj_5050, n9_adj_5051, 
        n9_adj_5052, n62, n12_adj_5053, n25796, n25797;
    wire [7:0]x_pl;   // g:/fpga/mxo2/system/project/oled12832.v(23[19:23])
    
    wire n25798, n23279, n23278, n23280, n8_adj_5054;
    wire [3:0]n4264;
    
    wire n14, n10_adj_5055, n25565, n15_adj_5056, n25789, n27, n26417, 
        n26495, n26497, n16743, n25646, n25763, n4_adj_5057, n26416, 
        n16320, n25764, n25713, n24, n25649, n9_adj_5058, n6028, 
        n25563, n26450, n25577, n25560, n26449, n26454, n23099, 
        n6_adj_5059, n7_adj_5060, n12_adj_5061, n25600, n25580, n23716, 
        n12_adj_5062, n26494, n23313, n25612, n25761, n12024, n23312, 
        n25678, n26493, n9_adj_5063, n25784, n24908, n25658, n25799, 
        n23674, n23345, n25620, n79, n6_adj_5064, n26, n25693, 
        n25760, n25497, n32_adj_5065, n25215, n25211, n25216;
    wire [4:0]n2535;
    
    wire n29_adj_5066, n26_adj_5067, n29_adj_5068, n32_adj_5069, n13581;
    wire [5:0]state_5__N_840;
    
    wire n25213, n25212, n25214, n25585, n25719, n25470, n23_adj_5070, 
        n23787, n21577, n25614, n25616, n18, n21575, n15_adj_5071, 
        n24914, n24915, n23590, n13, n24139, n25640, n2557, n23175, 
        n25684, clk_c_enable_1401, n16443, n5_adj_5072;
    wire [15:0]n141;
    wire [15:0]n167;
    
    wire n23507, n30, n11_adj_5073, n25788, n19, n16_adj_5074, n6_adj_5075, 
        n25036, n6550, n23229, n25581;
    wire [7:0]x_pl_7__N_529;
    wire [7:0]n3624;
    
    wire clk_c_enable_694;
    wire [7:0]n3536;
    
    wire n25191;
    wire [7:0]char_7__N_553;
    
    wire n25743, n43_adj_5076, n27_adj_5077, n6178, n20729, n24714, 
        n24713, n24715, n25745, n23153, n25750, n25749, n4_adj_5078, 
        n12_adj_5079, n22465, n25744, n5_adj_5080, n26455, n23350, 
        n23898, n25691, n25636, n25692, n4_adj_5081, n25074, n23769, 
        n23930, n23931, n23932, n23907, n25787, n23920, n23897, 
        n18_adj_5082, n22, n23895, n24711, n24710, n24712, n23867, 
        n23913, n23914, n25771, n26778, n23892, n25752, n25624, 
        n25791, n25790, n23755, n23941, n23906, n4_adj_5083, n25608, 
        clk_c_enable_1421, n24696, n24695, n24697, n25189, n20727, 
        n25121, n23_adj_5084, n16_adj_5085, n23927, n23928, n23929, 
        n23904, n23923, n23900, n24966, n25594, n25667, n7109, 
        n25872, n21029, n6_adj_5086, n23917, n4_adj_5087, n23894, 
        n24964, n24683, n23911, n23891, n6_adj_5088, n20788, n83, 
        n25756, n89, n58, n6_adj_5089, n23926, n23903;
    wire [15:0]cnt_c;   // g:/fpga/mxo2/system/project/oled12832.v(28[36:39])
    
    wire n20, n16_adj_5090, n25660, n8418, n16_adj_5091, n19_adj_5092, 
        n25186, n25187;
    wire [7:0]x_pl_7__N_700;
    
    wire n25578, n15856, n18_adj_5093, n25115, n4_adj_5094, clk_c_enable_1423, 
        n20715, n23718, n3264, n10049, n25683, n25769, n25770, 
        n16_adj_5095, n4_adj_5096, n25631, n8723, n16_adj_5097, n5_adj_5098, 
        n25674, n20_adj_5099, n25073, n15942, n25564, n25575, n23349, 
        n23589, n23803, n17773, n86, n25758, n23159, n60, n23157, 
        n62_adj_5100, n25694;
    wire [7:0]num1_7__N_724;
    
    wire n16391, n23869, n16678, n24049, n4432, n25609, clk_c_enable_1427, 
        n6_adj_5101, n25711, n25718, n25657, n25593, n23342;
    wire [7:0]char_reg_7__N_772;
    
    wire n25539, n25759, n20504, n20592, n23223, n20_adj_5102, n25677, 
        n4_adj_5103, n20591, n20590, n20503, n20502, n9817, n25639, 
        n20589, n20588, n25031, n20587, n25030, n4_adj_5104, n16_adj_5105, 
        n28, n31_adj_5106, n39;
    wire [7:0]char_7__N_756;
    
    wire n16111, n4_adj_5107, n23698, n8725, n20586, n16722, n25589, 
        n23942, n25123, n25122, n25124, n12017, n16_adj_5108, n24961, 
        n23945, n23761, n23946, n25119, n25590, n65, n41_adj_5109, 
        n24682, n24681, n20585, n16664, clk_c_enable_1436, n12019, 
        n20501;
    wire [1:0]n5817;
    
    wire n25034, n25035, n25605, n25622, n16_adj_5110, n25604, n25062, 
        n15_adj_5111, n15_adj_5112, n23958, n4_adj_5113, n24047, clk_c_enable_1429, 
        n20500, n68_adj_5114, n25579, n23306, n23307, n4_adj_5115, 
        n4434, n4_adj_5116;
    wire [0:0]n3189;
    
    wire n16_adj_5117, n74, n89_adj_5118, n20499, n76, n136, n20498, 
        n14_adj_5119, n15_adj_5120, n96, n105, n25044, n25047, n25048, 
        n23954, n16_adj_5121, n12116, n25570, n16_adj_5122, n93, 
        n25063, n16_adj_5123, n21240, n16_adj_5124, n37_adj_5125, 
        n25805, n61, n45, n4_adj_5126, n25046, n25045, n16_adj_5127, 
        n16_adj_5128, n25064, n20497, n23360, n24905, n11_adj_5129, 
        n21243, n16_adj_5130, n25037, n25412, n11_adj_5131, n16_adj_5132, 
        n27_adj_5133;
    wire [15:0]num1_delay_15__N_780;
    
    wire n25559, n16726, n23209, n15_adj_5134, n16_adj_5135, n16_adj_5136, 
        n25060, n16_adj_5137, n16_adj_5138, n8_adj_5139, n16_adj_5140;
    wire [63:0]n2030;
    wire [63:0]n2162;
    
    wire n25068, n20748, n25645, n23861, n16_adj_5141, n16_adj_5142, 
        n25672, n15_adj_5143, n16_adj_5144, n16_adj_5145, n25033, 
        n25032, n16_adj_5146, n16_adj_5147, n4_adj_5148, n16_adj_5149, 
        n16_adj_5150, n26451, n26453, n16_adj_5151, n16_adj_5152, 
        n9753, n35, n31_adj_5153;
    wire [5:0]state_back_5__N_858;
    
    wire n25653, n24_adj_5154, n25695, n25754, n42_adj_5155, n24_adj_5156, 
        n24_adj_5157, n24_adj_5158, n24_adj_5159, n94, n24_adj_5160, 
        n23318, n4_adj_5161, n25697, n25698, n24_adj_5162, n24_adj_5163, 
        n14_adj_5164, n10_adj_5165, n25665, n26777, n26042, n25762, 
        n25786, n24963, n24962, n11_adj_5166, n26039, n30_adj_5167, 
        n23821, n18_adj_5168, n50, n24187, n44, n20_adj_5169, n25496, 
        n22_adj_5170, n23935, n25748, n6170, n20573, n25671, n20572, 
        n20442, n20496, n25629, n17_adj_5171, n24_adj_5172, n20571, 
        n20495;
    wire [4:0]n331;
    
    wire n69_adj_5173, n13_adj_5174, n23947, n24906, n24907, n25324, 
        n20494, n20493, n20492, n23909, n23910, n23956, n23959, 
        n23915, n23916, n23918, n23919, n25556, n19_adj_5175, n6_adj_5176, 
        n21246, n19_adj_5177, n6_adj_5178, n20491, n25628, n13577, 
        n7110, n7112, n23314, n19_adj_5179, n6_adj_5180, n25310, 
        n20490, n20489, n23957, n25666, n23955, n5995, n9_adj_5181, 
        n8724, n17_adj_5182, n23310, n25641, n23921, n23922, n23924, 
        n23925, n6104, n25411, n8_adj_5183, n25598, n34_adj_5184, 
        n23965, n23504, n23378, n23359, n23939, n23940, n72, n23379;
    wire [7:0]n361;
    
    wire n14_adj_5185, n23963, n23964, n25428, n7_adj_5186, n25804, 
        n25871, n25810, n25809, n25803, n25430, n20526, n20525, 
        n23878, n8876, n20524, n20523, n25821, n25822, n25427, 
        n25431, n25429, n20522, n20521, n20520, n20519, n25410;
    
    LUT4 state_5__I_0_377_i11_2_lut_rep_355_3_lut_4_lut (.A(state[5]), .B(state[4]), 
         .C(n8), .D(state[3]), .Z(n25637)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam state_5__I_0_377_i11_2_lut_rep_355_3_lut_4_lut.init = 16'hfffe;
    LUT4 i21000_3_lut (.A(char_reg[6]), .B(char_reg[2]), .C(cnt_write[3]), 
         .Z(n23877)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21000_3_lut.init = 16'hcaca;
    LUT4 i17793_3_lut_4_lut (.A(n25635), .B(n25630), .C(n23422), .D(n25601), 
         .Z(n17)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(139[72:96])
    defparam i17793_3_lut_4_lut.init = 16'h0001;
    PFUMX i66 (.BLUT(n32), .ALUT(n37), .C0(cnt_main[3]), .Z(n43));
    FD1P3IX cnt_delay_i0_i4 (.D(n2559[4]), .SP(clk_c_enable_1452), .CD(n12055), 
            .CK(clk_c), .Q(cnt_delay[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam cnt_delay_i0_i4.GSR = "ENABLED";
    FD1P3AX cnt_init_i0_i0 (.D(n3871[0]), .SP(clk_c_enable_1359), .CK(clk_c), 
            .Q(cnt_init[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam cnt_init_i0_i0.GSR = "ENABLED";
    FD1P3AY y_ph_i0_i0 (.D(n5820[0]), .SP(clk_c_enable_690), .CK(clk_c), 
            .Q(y_ph[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam y_ph_i0_i0.GSR = "ENABLED";
    FD1P3AX char_reg_i0_i0 (.D(n3492[0]), .SP(clk_c_enable_702), .CK(clk_c), 
            .Q(char_reg[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam char_reg_i0_i0.GSR = "ENABLED";
    FD1S3AY num1_delay_i0 (.D(num1_delay_15__N_605[0]), .CK(clk_c), .Q(num1_delay[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam num1_delay_i0.GSR = "ENABLED";
    FD1S3AY state_back_i0 (.D(state_back_5__N_659[0]), .CK(clk_c), .Q(state_back[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam state_back_i0.GSR = "ENABLED";
    FD1P3AY oled_csn_368 (.D(n3153[0]), .SP(clk_c_enable_10), .CK(clk_c), 
            .Q(oled_csn_c)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam oled_csn_368.GSR = "ENABLED";
    LUT4 i2651_2_lut_3_lut (.A(cnt_init[0]), .B(cnt_init[1]), .C(cnt_init[2]), 
         .Z(n1[2])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(41[4] 175[11])
    defparam i2651_2_lut_3_lut.init = 16'h7878;
    FD1S3AY x_ph_i0 (.D(x_ph_7__N_519[0]), .CK(clk_c), .Q(x_ph[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam x_ph_i0.GSR = "ENABLED";
    LUT4 i21489_2_lut_3_lut_4_lut (.A(n9), .B(n25587), .C(clk_c_enable_1352), 
         .D(n16632), .Z(clk_c_enable_114)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (C)) */ ;
    defparam i21489_2_lut_3_lut_4_lut.init = 16'hd0f0;
    L6MUX21 i22037 (.D0(n25374), .D1(n25371), .SD(n25574), .Z(n23953));
    LUT4 i21421_2_lut_3_lut_4_lut (.A(n9), .B(n25587), .C(clk_c_enable_1352), 
         .D(n16666), .Z(clk_c_enable_690)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (C)) */ ;
    defparam i21421_2_lut_3_lut_4_lut.init = 16'hd0f0;
    PFUMX i22035 (.BLUT(n25373), .ALUT(n25372), .C0(n25635), .Z(n25374));
    LUT4 i3_4_lut (.A(state[1]), .B(n36), .C(n25610), .D(state[2]), 
         .Z(n5)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(41[4] 175[11])
    defparam i3_4_lut.init = 16'h0020;
    PFUMX i22032 (.BLUT(n25561), .ALUT(n25369), .C0(cnt_scan[0]), .Z(n25371));
    PFUMX i34 (.BLUT(n16), .ALUT(n20791), .C0(cnt_scan[3]), .Z(n3599));
    LUT4 i20999_3_lut (.A(char_reg[5]), .B(char_reg[1]), .C(cnt_write[3]), 
         .Z(n23876)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20999_3_lut.init = 16'hcaca;
    LUT4 i20998_3_lut (.A(char_reg[7]), .B(char_reg[3]), .C(cnt_write[3]), 
         .Z(n23875)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20998_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_rep_287 (.A(n29), .B(state[3]), .C(n16393), .D(n9173), 
         .Z(clk_c_enable_1431)) /* synthesis lut_function=(A (B (C (D))+!B (C))) */ ;
    defparam i1_4_lut_rep_287.init = 16'ha020;
    FD1P3IX cnt_delay_i0_i3 (.D(n2559[3]), .SP(clk_c_enable_1452), .CD(n12055), 
            .CK(clk_c), .Q(cnt_delay[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam cnt_delay_i0_i3.GSR = "ENABLED";
    FD1P3IX cnt_delay_i0_i2 (.D(n2559[2]), .SP(clk_c_enable_1452), .CD(n12055), 
            .CK(clk_c), .Q(cnt_delay[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam cnt_delay_i0_i2.GSR = "ENABLED";
    FD1P3IX cnt_delay_i0_i1 (.D(n2559[1]), .SP(clk_c_enable_1452), .CD(n12055), 
            .CK(clk_c), .Q(cnt_delay[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam cnt_delay_i0_i1.GSR = "ENABLED";
    FD1P3IX num2_i0_i7 (.D(num2_7__N_748[7]), .SP(clk_c_enable_1431), .CD(n12049), 
            .CK(clk_c), .Q(num2[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam num2_i0_i7.GSR = "ENABLED";
    FD1P3IX num2_i0_i6 (.D(num2_7__N_748[6]), .SP(clk_c_enable_1431), .CD(n12049), 
            .CK(clk_c), .Q(num2[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam num2_i0_i6.GSR = "ENABLED";
    FD1P3IX num2_i0_i5 (.D(num2_7__N_748[5]), .SP(clk_c_enable_1431), .CD(n12049), 
            .CK(clk_c), .Q(num2[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam num2_i0_i5.GSR = "ENABLED";
    FD1P3IX num2_i0_i4 (.D(num2_7__N_748[4]), .SP(clk_c_enable_1431), .CD(n12049), 
            .CK(clk_c), .Q(num2[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam num2_i0_i4.GSR = "ENABLED";
    FD1P3IX num2_i0_i3 (.D(num2_7__N_748[3]), .SP(clk_c_enable_1431), .CD(n12049), 
            .CK(clk_c), .Q(num2[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam num2_i0_i3.GSR = "ENABLED";
    FD1P3IX num2_i0_i2 (.D(num2_7__N_748[2]), .SP(clk_c_enable_1431), .CD(n12049), 
            .CK(clk_c), .Q(num2[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam num2_i0_i2.GSR = "ENABLED";
    FD1P3IX num1_i0_i4 (.D(num1_7__N_732[4]), .SP(clk_c_enable_1432), .CD(n14556), 
            .CK(clk_c), .Q(num1[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam num1_i0_i4.GSR = "ENABLED";
    FD1P3IX num1_i0_i2 (.D(num1_7__N_732[2]), .SP(clk_c_enable_1432), .CD(n14556), 
            .CK(clk_c), .Q(num1[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam num1_i0_i2.GSR = "ENABLED";
    FD1P3IX num1_i0_i1 (.D(num1_7__N_732[1]), .SP(clk_c_enable_1432), .CD(n14556), 
            .CK(clk_c), .Q(num1[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam num1_i0_i1.GSR = "ENABLED";
    FD1P3AX y_pl_i0_i1 (.D(n16636), .SP(clk_c_enable_114), .CK(clk_c), 
            .Q(y_pl[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam y_pl_i0_i1.GSR = "ENABLED";
    FD1P3IX cnt_scan_i0_i0 (.D(cnt_scan_4__N_682[0]), .SP(clk_c_enable_1446), 
            .CD(n12042), .CK(clk_c), .Q(cnt_scan[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam cnt_scan_i0_i0.GSR = "ENABLED";
    FD1P3IX cnt_main_1988__i0 (.D(n2[0]), .SP(clk_c_enable_1352), .CD(n12039), 
            .CK(clk_c), .Q(cnt_main[0]));   // g:/fpga/mxo2/system/project/oled12832.v(53[12:40])
    defparam cnt_main_1988__i0.GSR = "ENABLED";
    LUT4 i9238_2_lut_3_lut (.A(n29), .B(state[3]), .C(n16393), .Z(n12049)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i9238_2_lut_3_lut.init = 16'h2020;
    LUT4 n25039_bdd_3_lut_4_lut (.A(n25808), .B(n25558), .C(state[3]), 
         .D(n25038), .Z(n25040)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;
    defparam n25039_bdd_3_lut_4_lut.init = 16'hf808;
    LUT4 i2_3_lut_rep_275 (.A(n23134), .B(n1358), .C(n1359), .Z(n25557)) /* synthesis lut_function=(A+(B+(C))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(129[51:75])
    defparam i2_3_lut_rep_275.init = 16'hfefe;
    LUT4 n9304_bdd_4_lut_22661 (.A(n9304), .B(n322), .C(cnt_scan[0]), 
         .D(cnt_scan[3]), .Z(n25469)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (B (C+!(D))+!B (C (D)+!C !(D)))) */ ;
    defparam n9304_bdd_4_lut_22661.init = 16'hf0c5;
    LUT4 i20868_2_lut_rep_279_3_lut_3_lut (.A(n25635), .B(num2[0]), .C(n25676), 
         .Z(n25561)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(111[7] 142[14])
    defparam i20868_2_lut_rep_279_3_lut_3_lut.init = 16'h4040;
    LUT4 i1_4_lut (.A(n15), .B(n25696), .C(n25823), .D(cnt_scan[4]), 
         .Z(n23311)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(41[4] 175[11])
    defparam i1_4_lut.init = 16'hc088;
    LUT4 i21259_3_lut (.A(n23311), .B(n21), .C(state[5]), .Z(n23)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(41[4] 175[11])
    defparam i21259_3_lut.init = 16'hcaca;
    PFUMX i101 (.BLUT(n9872), .ALUT(n20744), .C0(cnt_main[2]), .Z(n59));
    LUT4 i13259_2_lut (.A(state[4]), .B(state_back[0]), .Z(n41)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i13259_2_lut.init = 16'h1111;
    LUT4 i1_4_lut_adj_73 (.A(state[4]), .B(state[0]), .C(n25682), .D(n25638), 
         .Z(n34)) /* synthesis lut_function=(!((B (C+!(D))+!B (C (D)))+!A)) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(41[4] 175[11])
    defparam i1_4_lut_adj_73.init = 16'h0a22;
    PFUMX i135 (.BLUT(n102), .ALUT(n80), .C0(cnt_main[2]), .Z(n99));
    LUT4 n2421_bdd_4_lut_21994_4_lut (.A(n25635), .B(n25676), .C(n25601), 
         .D(n23763), .Z(n25311)) /* synthesis lut_function=(!(A ((D)+!C)+!A !(B))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(111[7] 142[14])
    defparam n2421_bdd_4_lut_21994_4_lut.init = 16'h44e4;
    LUT4 i20726_2_lut_3_lut_4_lut (.A(n25651), .B(oled_dcn_N_888), .C(state_back[5]), 
         .D(n25755), .Z(n23579)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;
    defparam i20726_2_lut_3_lut_4_lut.init = 16'hf080;
    LUT4 i20727_2_lut_3_lut_4_lut (.A(n25651), .B(oled_dcn_N_888), .C(state_back[4]), 
         .D(n25755), .Z(n23581)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;
    defparam i20727_2_lut_3_lut_4_lut.init = 16'hf080;
    LUT4 i20728_2_lut_3_lut_4_lut (.A(n25651), .B(oled_dcn_N_888), .C(state_back[0]), 
         .D(n25755), .Z(n23583)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;
    defparam i20728_2_lut_3_lut_4_lut.init = 16'hf080;
    LUT4 n23706_bdd_3_lut_4_lut_4_lut (.A(n25635), .B(n25601), .C(n25676), 
         .D(n25753), .Z(n25120)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A !(B (C (D))))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(111[7] 142[14])
    defparam n23706_bdd_3_lut_4_lut_4_lut.init = 16'h4080;
    LUT4 n2533_bdd_2_lut (.A(state_back[5]), .B(state[4]), .Z(n25495)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam n2533_bdd_2_lut.init = 16'h2222;
    LUT4 i6048_4_lut_4_lut_4_lut_4_lut_4_lut (.A(n25635), .B(n25753), .C(n25601), 
         .D(n25676), .Z(n8855)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A !(B (C (D)+!C !(D))+!B !(C+(D))))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(111[7] 142[14])
    defparam i6048_4_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h6a0f;
    LUT4 mux_131_Mux_7_i12_3_lut (.A(n1138), .B(n1278), .C(cnt_scan[0]), 
         .Z(n12)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(111[7] 142[14])
    defparam mux_131_Mux_7_i12_3_lut.init = 16'hcaca;
    LUT4 i13524_2_lut (.A(n998), .B(cnt_scan[0]), .Z(n11)) /* synthesis lut_function=(A (B)) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(111[7] 142[14])
    defparam i13524_2_lut.init = 16'h8888;
    LUT4 mux_131_Mux_6_i9_3_lut (.A(n579), .B(n719), .C(cnt_scan[0]), 
         .Z(n9_adj_5037)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(111[7] 142[14])
    defparam mux_131_Mux_6_i9_3_lut.init = 16'hcaca;
    LUT4 i13526_2_lut (.A(n439), .B(cnt_scan[0]), .Z(n8_adj_5038)) /* synthesis lut_function=(A (B)) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(111[7] 142[14])
    defparam i13526_2_lut.init = 16'h8888;
    PFUMX i22174 (.BLUT(n25800), .ALUT(n25801), .C0(cnt_main[1]), .Z(n9));
    LUT4 mux_131_Mux_7_i9_3_lut (.A(n578), .B(n718), .C(cnt_scan[0]), 
         .Z(n9_adj_5039)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(111[7] 142[14])
    defparam mux_131_Mux_7_i9_3_lut.init = 16'hcaca;
    LUT4 i13523_2_lut (.A(n438), .B(cnt_scan[0]), .Z(n8_adj_5040)) /* synthesis lut_function=(A (B)) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(111[7] 142[14])
    defparam i13523_2_lut.init = 16'h8888;
    LUT4 i13364_3_lut (.A(n1357), .B(n23415), .C(n1356), .Z(n31)) /* synthesis lut_function=(!(A (B+!(C))+!A (B+(C)))) */ ;
    defparam i13364_3_lut.init = 16'h2121;
    PFUMX i22001 (.BLUT(n25325), .ALUT(n25323), .C0(state[3]), .Z(n25326));
    LUT4 n23966_bdd_4_lut (.A(n23966), .B(n23967), .C(cnt[4]), .D(n25558), 
         .Z(n25553)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam n23966_bdd_4_lut.init = 16'hca00;
    LUT4 n9339_bdd_4_lut_22150 (.A(n25686), .B(state[4]), .C(cnt_scan[3]), 
         .D(cnt_scan[0]), .Z(n25519)) /* synthesis lut_function=(!(A (C)+!A !(B+(C+!(D))))) */ ;
    defparam n9339_bdd_4_lut_22150.init = 16'h5e5f;
    LUT4 i1_4_lut_adj_74 (.A(cnt_init[0]), .B(num1_delay[0]), .C(n15_adj_5041), 
         .D(n25650), .Z(n23253)) /* synthesis lut_function=(!(A (B (D))+!A (B (C+(D))+!B (C)))) */ ;
    defparam i1_4_lut_adj_74.init = 16'h23af;
    LUT4 mux_131_Mux_4_i12_3_lut (.A(n1141), .B(n1281), .C(cnt_scan[0]), 
         .Z(n12_adj_5042)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(111[7] 142[14])
    defparam mux_131_Mux_4_i12_3_lut.init = 16'hcaca;
    LUT4 i13217_4_lut (.A(n25599), .B(n25566), .C(n92), .D(cnt_scan[0]), 
         .Z(n10074)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(111[7] 142[14])
    defparam i13217_4_lut.init = 16'hc088;
    PFUMX i21997 (.BLUT(n25315), .ALUT(n25314), .C0(cnt_scan[1]), .Z(n25316));
    LUT4 mux_131_Mux_5_i12_3_lut (.A(n1140), .B(n1280), .C(cnt_scan[0]), 
         .Z(n12_adj_5043)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(111[7] 142[14])
    defparam mux_131_Mux_5_i12_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_75 (.A(n25566), .B(n25599), .C(n25621), .D(cnt_scan[0]), 
         .Z(n22121)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(111[7] 142[14])
    defparam i1_4_lut_adj_75.init = 16'ha088;
    LUT4 i17809_2_lut_3_lut_4_lut_4_lut (.A(n25635), .B(n25601), .C(n23422), 
         .D(n25630), .Z(n17_adj_5044)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(111[7] 142[14])
    defparam i17809_2_lut_3_lut_4_lut_4_lut.init = 16'h0008;
    FD1P3AY state_i0_i0 (.D(n42), .SP(clk_c_enable_1374), .CK(clk_c), 
            .Q(state[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam state_i0_i0.GSR = "ENABLED";
    LUT4 i69_4_lut (.A(cnt_main[0]), .B(time_data[5]), .C(cnt_main[1]), 
         .D(\tamp_data[1] ), .Z(n46)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C)) */ ;
    defparam i69_4_lut.init = 16'h8f85;
    LUT4 i1_4_lut_adj_76 (.A(cnt_scan[2]), .B(x_ph[0]), .C(n865), .D(cnt_scan[3]), 
         .Z(n12_adj_5045)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam i1_4_lut_adj_76.init = 16'ha088;
    PFUMX i21995 (.BLUT(n25312), .ALUT(n25311), .C0(n25574), .Z(n25313));
    LUT4 cnt_3__bdd_3_lut_22139 (.A(cnt[0]), .B(cnt[4]), .C(cnt[1]), .Z(n25537)) /* synthesis lut_function=(!(A+(B (C)))) */ ;
    defparam cnt_3__bdd_3_lut_22139.init = 16'h1515;
    LUT4 i20830_3_lut_4_lut_4_lut (.A(n25635), .B(n25753), .C(n25676), 
         .D(n25601), .Z(n23694)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(111[7] 142[14])
    defparam i20830_3_lut_4_lut_4_lut.init = 16'h4000;
    LUT4 i1_2_lut_3_lut (.A(state[2]), .B(n25586), .C(state_back[5]), 
         .Z(n23281)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h1010;
    LUT4 i2_3_lut_4_lut_4_lut (.A(n25635), .B(n23347), .C(n25601), .D(n25632), 
         .Z(n23348)) /* synthesis lut_function=(A (B (C (D)))+!A !(((D)+!C)+!B)) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(111[7] 142[14])
    defparam i2_3_lut_4_lut_4_lut.init = 16'h8040;
    LUT4 cnt_3__bdd_3_lut (.A(cnt[0]), .B(cnt[2]), .C(cnt[1]), .Z(n25538)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)+!B !(C)))) */ ;
    defparam cnt_3__bdd_3_lut.init = 16'h4949;
    LUT4 mux_131_Mux_3_i9_3_lut (.A(n582), .B(n722), .C(cnt_scan[0]), 
         .Z(n9_adj_5046)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(111[7] 142[14])
    defparam mux_131_Mux_3_i9_3_lut.init = 16'hcaca;
    LUT4 time_data_0__bdd_4_lut_then_4_lut (.A(char[1]), .B(cnt_main[2]), 
         .C(cnt_main[3]), .D(cnt_main[4]), .Z(n25785)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam time_data_0__bdd_4_lut_then_4_lut.init = 16'h02c2;
    LUT4 mux_131_Mux_4_i9_3_lut (.A(n581), .B(n721), .C(cnt_scan[0]), 
         .Z(n9_adj_5047)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(111[7] 142[14])
    defparam mux_131_Mux_4_i9_3_lut.init = 16'hcaca;
    PFUMX i15043 (.BLUT(n68), .ALUT(n69), .C0(cnt_scan[2]), .Z(n7));
    PFUMX mux_131_Mux_1_i6 (.BLUT(n4), .ALUT(n5_adj_5048), .C0(cnt_scan[1]), 
          .Z(n6)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;
    L6MUX21 i21004 (.D0(n23879), .D1(n23880), .SD(cnt_write[1]), .Z(n23881));
    LUT4 mux_131_Mux_6_i12_3_lut (.A(n1139), .B(n1279), .C(cnt_scan[0]), 
         .Z(n12_adj_5049)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(111[7] 142[14])
    defparam mux_131_Mux_6_i12_3_lut.init = 16'hcaca;
    LUT4 mux_131_Mux_6_i11_4_lut (.A(n23134), .B(n999), .C(cnt_scan[0]), 
         .D(n23415), .Z(n11_adj_5050)) /* synthesis lut_function=(A (B (C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(111[7] 142[14])
    defparam mux_131_Mux_6_i11_4_lut.init = 16'hc0c5;
    LUT4 mux_131_Mux_2_i9_3_lut (.A(n583), .B(n723), .C(cnt_scan[0]), 
         .Z(n9_adj_5051)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(111[7] 142[14])
    defparam mux_131_Mux_2_i9_3_lut.init = 16'hcaca;
    LUT4 mux_131_Mux_5_i9_3_lut (.A(n580), .B(n720), .C(cnt_scan[0]), 
         .Z(n9_adj_5052)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(111[7] 142[14])
    defparam mux_131_Mux_5_i9_3_lut.init = 16'hcaca;
    LUT4 mux_415_Mux_29_i62_4_lut (.A(n25599), .B(n23415), .C(n1356), 
         .D(n1357), .Z(n62)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)+!C !(D)))+!A (B+((D)+!C)))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(129[51:75])
    defparam mux_415_Mux_29_i62_4_lut.init = 16'h0a30;
    LUT4 mux_131_Mux_3_i12_3_lut (.A(n1142), .B(n1282), .C(cnt_scan[0]), 
         .Z(n12_adj_5053)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(111[7] 142[14])
    defparam mux_131_Mux_3_i12_3_lut.init = 16'hcaca;
    PFUMX i22171 (.BLUT(n25796), .ALUT(n25797), .C0(x_pl[4]), .Z(n25798));
    LUT4 i1_2_lut_3_lut_adj_77 (.A(state[2]), .B(n25586), .C(state_back[4]), 
         .Z(n23279)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_77.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_78 (.A(state[2]), .B(n25586), .C(state_back[0]), 
         .Z(n23278)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_78.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_79 (.A(state[2]), .B(n25586), .C(state_back[2]), 
         .Z(n23280)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_79.init = 16'h1010;
    LUT4 i2_3_lut_rep_319 (.A(num2[4]), .B(char[4]), .C(n8_adj_5054), 
         .Z(n25601)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;
    defparam i2_3_lut_rep_319.init = 16'h9696;
    LUT4 mux_1622_i2_4_lut (.A(n9304), .B(n322), .C(cnt_scan[3]), .D(cnt_scan[0]), 
         .Z(n4264[1])) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+(D))+!B !(C (D)+!C !(D))))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(101[30] 110[58])
    defparam mux_1622_i2_4_lut.init = 16'h3005;
    LUT4 i7_4_lut (.A(num1[0]), .B(n14), .C(n10_adj_5055), .D(num1[6]), 
         .Z(n9304)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(102[11:15])
    defparam i7_4_lut.init = 16'hfffe;
    LUT4 i6_4_lut (.A(num1[3]), .B(num1[1]), .C(num1[5]), .D(num1[7]), 
         .Z(n14)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(102[11:15])
    defparam i6_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut (.A(num1[2]), .B(num1[4]), .Z(n10_adj_5055)) /* synthesis lut_function=(A+(B)) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(102[11:15])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i21564_2_lut_rep_283_2_lut_4_lut (.A(num2[4]), .B(char[4]), .C(n8_adj_5054), 
         .D(n25635), .Z(n25565)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C+(D)))+!A (B (C+(D))+!B ((D)+!C))) */ ;
    defparam i21564_2_lut_rep_283_2_lut_4_lut.init = 16'hff69;
    LUT4 i18105_1_lut_rep_292_3_lut (.A(num2[4]), .B(char[4]), .C(n8_adj_5054), 
         .Z(n25574)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B (C)+!B !(C)))) */ ;
    defparam i18105_1_lut_rep_292_3_lut.init = 16'h6969;
    LUT4 i13261_4_lut (.A(state[2]), .B(n15_adj_5056), .C(n25789), .D(cnt_scan[4]), 
         .Z(n27)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B (C (D))))) */ ;
    defparam i13261_4_lut.init = 16'h0511;
    LUT4 n25601_bdd_3_lut_22514 (.A(n25635), .B(n25676), .C(cnt_scan[0]), 
         .Z(n26417)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;
    defparam n25601_bdd_3_lut_22514.init = 16'h0404;
    LUT4 n26496_bdd_2_lut_3_lut (.A(n26495), .B(state[4]), .C(state[1]), 
         .Z(n26497)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;
    defparam n26496_bdd_2_lut_3_lut.init = 16'h0202;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut (.A(cnt_main[1]), .B(n16743), .C(n25646), 
         .D(n25763), .Z(n4_adj_5057)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A ((C)+!B))) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut.init = 16'h0c04;
    LUT4 n25601_bdd_4_lut_22515 (.A(n25635), .B(n25676), .C(n25753), .D(cnt_scan[0]), 
         .Z(n26416)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(D)))) */ ;
    defparam n25601_bdd_4_lut_22515.init = 16'h60f7;
    LUT4 i13543_2_lut_2_lut_4_lut (.A(num2[4]), .B(char[4]), .C(n8_adj_5054), 
         .D(cnt_scan[0]), .Z(n16320)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C+(D)))+!A (B (C+(D))+!B ((D)+!C))) */ ;
    defparam i13543_2_lut_2_lut_4_lut.init = 16'hff69;
    LUT4 i1_4_lut_adj_80 (.A(num1_delay[0]), .B(n25755), .C(n25651), .D(oled_dcn_N_888), 
         .Z(n15_adj_5041)) /* synthesis lut_function=(A (B+(C))+!A !((D)+!C)) */ ;
    defparam i1_4_lut_adj_80.init = 16'ha8f8;
    LUT4 i13615_2_lut_4_lut (.A(cnt_main[4]), .B(n25764), .C(cnt_main[3]), 
         .D(n25713), .Z(n16393)) /* synthesis lut_function=(A (D)+!A (B ((D)+!C)+!B (C+(D)))) */ ;
    defparam i13615_2_lut_4_lut.init = 16'hff14;
    LUT4 i1_4_lut_adj_81 (.A(n24), .B(state_back[0]), .C(n25649), .D(n9_adj_5058), 
         .Z(state_back_5__N_659[0])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A ((D)+!B))) */ ;
    defparam i1_4_lut_adj_81.init = 16'h0ace;
    LUT4 cnt_scan_2__bdd_4_lut_22558 (.A(n25601), .B(num2[0]), .C(n6028), 
         .D(n25563), .Z(n26450)) /* synthesis lut_function=(!(A (B+(C))+!A (B+!(D)))) */ ;
    defparam cnt_scan_2__bdd_4_lut_22558.init = 16'h1302;
    LUT4 cnt_scan_2__bdd_4_lut_22521 (.A(n25601), .B(n25577), .C(n25560), 
         .D(num2[0]), .Z(n26449)) /* synthesis lut_function=(!(A (B+(D))+!A !(C))) */ ;
    defparam cnt_scan_2__bdd_4_lut_22521.init = 16'h5072;
    LUT4 i1_2_lut_3_lut_4_lut (.A(cnt_scan[0]), .B(n25686), .C(cnt_scan[4]), 
         .D(cnt_scan[3]), .Z(n9173)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0020;
    LUT4 n1424_bdd_3_lut (.A(n1424), .B(cnt_scan[2]), .C(cnt_scan[1]), 
         .Z(n26454)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;
    defparam n1424_bdd_3_lut.init = 16'h0202;
    PFUMX mux_131_Mux_5_i7 (.BLUT(n23099), .ALUT(n6_adj_5059), .C0(cnt_scan[2]), 
          .Z(n7_adj_5060)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;
    LUT4 mux_131_Mux_1_i12_3_lut (.A(n1144), .B(n1284), .C(cnt_scan[0]), 
         .Z(n12_adj_5061)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(111[7] 142[14])
    defparam mux_131_Mux_1_i12_3_lut.init = 16'hcaca;
    LUT4 i3208_3_lut_4_lut_4_lut (.A(n25600), .B(n25580), .C(n25601), 
         .D(n25635), .Z(n23716)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A !(B+(C)))) */ ;
    defparam i3208_3_lut_4_lut_4_lut.init = 16'h5cfc;
    LUT4 mux_131_Mux_2_i12_3_lut (.A(n1143), .B(n1283), .C(cnt_scan[0]), 
         .Z(n12_adj_5062)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(111[7] 142[14])
    defparam mux_131_Mux_2_i12_3_lut.init = 16'hcaca;
    LUT4 n26494_bdd_3_lut (.A(n26494), .B(n23), .C(state[3]), .Z(n26495)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n26494_bdd_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_82 (.A(n23313), .B(n25612), .C(n25761), .D(n8), 
         .Z(n12024)) /* synthesis lut_function=(A (B)+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_82.init = 16'hc888;
    LUT4 i2_4_lut (.A(n23312), .B(state[0]), .C(n25678), .D(cnt_init[0]), 
         .Z(n23313)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i2_4_lut.init = 16'h0200;
    LUT4 i2644_2_lut (.A(cnt_init[1]), .B(cnt_init[0]), .Z(n1[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(79[49:64])
    defparam i2644_2_lut.init = 16'h6666;
    LUT4 i1_2_lut (.A(state[2]), .B(state[1]), .Z(n23312)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut.init = 16'h2222;
    LUT4 n25651_bdd_4_lut (.A(n25651), .B(state[0]), .C(state[2]), .D(cnt_init[0]), 
         .Z(n26493)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)))+!A ((C)+!B))) */ ;
    defparam n25651_bdd_4_lut.init = 16'h2c0c;
    LUT4 mux_131_Mux_1_i9_3_lut (.A(n584), .B(n724), .C(cnt_scan[0]), 
         .Z(n9_adj_5063)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(111[7] 142[14])
    defparam mux_131_Mux_1_i9_3_lut.init = 16'hcaca;
    LUT4 time_data_0__bdd_4_lut_else_4_lut (.A(char[1]), .B(cnt_main[2]), 
         .C(cnt_main[3]), .Z(n25784)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;
    defparam time_data_0__bdd_4_lut_else_4_lut.init = 16'h0202;
    LUT4 n23412_bdd_4_lut_21946 (.A(n25686), .B(cnt_scan[0]), .C(cnt_scan[3]), 
         .D(cnt_scan[4]), .Z(n24908)) /* synthesis lut_function=(!(A (C)+!A !(B (C+!(D))+!B ((D)+!C)))) */ ;
    defparam n23412_bdd_4_lut_21946.init = 16'h5b4f;
    LUT4 cnt_main_3__bdd_4_lut_22218 (.A(cnt_main[3]), .B(n25658), .C(cnt_main[1]), 
         .D(cnt_main[0]), .Z(n25799)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (C (D)+!C !(D)))) */ ;
    defparam cnt_main_3__bdd_4_lut_22218.init = 16'h0fd0;
    LUT4 i1_2_lut_adj_83 (.A(state[5]), .B(n23674), .Z(n23345)) /* synthesis lut_function=(!((B)+!A)) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(41[4] 175[11])
    defparam i1_2_lut_adj_83.init = 16'h2222;
    LUT4 i1_4_lut_adj_84 (.A(state[2]), .B(state[5]), .C(n25620), .D(n79), 
         .Z(n6_adj_5064)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(41[4] 175[11])
    defparam i1_4_lut_adj_84.init = 16'ha0a8;
    LUT4 i1_4_lut_adj_85 (.A(n26), .B(n25693), .C(n25760), .D(n25497), 
         .Z(n32_adj_5065)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B+!(D)))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(41[4] 175[11])
    defparam i1_4_lut_adj_85.init = 16'h3b0a;
    PFUMX i21941 (.BLUT(n25215), .ALUT(n25211), .C0(cnt_scan[1]), .Z(n25216));
    LUT4 i2716_2_lut (.A(cnt_write[1]), .B(cnt_write[0]), .Z(n2535[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(146[25:41])
    defparam i2716_2_lut.init = 16'h6666;
    LUT4 i13845_3_lut_4_lut (.A(cnt_scan[0]), .B(n25686), .C(n23694), 
         .D(num2[0]), .Z(n29_adj_5066)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(111[7] 142[14])
    defparam i13845_3_lut_4_lut.init = 16'h1000;
    LUT4 i13379_2_lut_3_lut_4_lut (.A(cnt_scan[0]), .B(n25686), .C(state[1]), 
         .D(cnt_scan[3]), .Z(n15)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(111[7] 142[14])
    defparam i13379_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i1_4_lut_adj_86 (.A(n26_adj_5067), .B(n29_adj_5068), .C(n25760), 
         .D(n25693), .Z(n32_adj_5069)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A ((D)+!B))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(41[4] 175[11])
    defparam i1_4_lut_adj_86.init = 16'h0ace;
    LUT4 i47_4_lut (.A(state[2]), .B(state[3]), .C(n13581), .D(state_5__N_840[4]), 
         .Z(n26_adj_5067)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(41[4] 175[11])
    defparam i47_4_lut.init = 16'h6420;
    PFUMX i21939 (.BLUT(n25213), .ALUT(n25212), .C0(n1355), .Z(n25214));
    LUT4 i1_2_lut_rep_303_3_lut_4_lut (.A(cnt_scan[0]), .B(n25686), .C(cnt_scan[4]), 
         .D(cnt_scan[3]), .Z(n25585)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(111[7] 142[14])
    defparam i1_2_lut_rep_303_3_lut_4_lut.init = 16'hfeff;
    LUT4 i13200_2_lut_3_lut_4_lut (.A(cnt_scan[0]), .B(n25686), .C(state[0]), 
         .D(cnt_scan[3]), .Z(n15_adj_5056)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(111[7] 142[14])
    defparam i13200_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 n9304_bdd_3_lut_4_lut (.A(cnt_scan[2]), .B(n25719), .C(cnt_scan[3]), 
         .D(cnt_scan[4]), .Z(n25470)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam n9304_bdd_3_lut_4_lut.init = 16'h7f80;
    LUT4 i1_4_lut_adj_87 (.A(state[4]), .B(n23_adj_5070), .C(n23787), 
         .D(state[3]), .Z(n21577)) /* synthesis lut_function=(!(A+(B (C (D))+!B (C+!(D))))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(41[4] 175[11])
    defparam i1_4_lut_adj_87.init = 16'h0544;
    LUT4 i20810_4_lut (.A(state[2]), .B(n25614), .C(n25616), .D(cnt_scan[4]), 
         .Z(n23674)) /* synthesis lut_function=(A+!(B (C (D))+!B (C+!(D)))) */ ;
    defparam i20810_4_lut.init = 16'hafee;
    LUT4 i2_3_lut (.A(n18), .B(state[3]), .C(state[4]), .Z(n21575)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(41[4] 175[11])
    defparam i2_3_lut.init = 16'h0202;
    LUT4 i31_4_lut (.A(n15_adj_5071), .B(state_back[2]), .C(state[5]), 
         .D(n25761), .Z(n18)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(41[4] 175[11])
    defparam i31_4_lut.init = 16'hca0a;
    LUT4 n24914_bdd_2_lut (.A(n24914), .B(cnt_main[4]), .Z(n24915)) /* synthesis lut_function=(A+(B)) */ ;
    defparam n24914_bdd_2_lut.init = 16'heeee;
    LUT4 i21424_4_lut (.A(state[1]), .B(n25637), .C(n23590), .D(n13), 
         .Z(n24139)) /* synthesis lut_function=(!(A+(B (C)+!B (C+(D))))) */ ;
    defparam i21424_4_lut.init = 16'h0405;
    LUT4 i13159_2_lut_rep_273_4_lut (.A(n25640), .B(state[4]), .C(state[5]), 
         .D(n2557), .Z(clk_c_enable_1374)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(169[5:10])
    defparam i13159_2_lut_rep_273_4_lut.init = 16'hffef;
    LUT4 i21378_4_lut (.A(n23175), .B(n25684), .C(n25761), .D(state[0]), 
         .Z(clk_c_enable_1401)) /* synthesis lut_function=(A+!(B+!(C (D)))) */ ;
    defparam i21378_4_lut.init = 16'hbaaa;
    LUT4 i3_4_lut_adj_88 (.A(cnt_init[0]), .B(n16443), .C(n5_adj_5072), 
         .D(n25651), .Z(n23175)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i3_4_lut_adj_88.init = 16'h1000;
    LUT4 i18_2_lut (.A(state[0]), .B(state[2]), .Z(n5_adj_5072)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(29[13:18])
    defparam i18_2_lut.init = 16'h6666;
    LUT4 i13720_2_lut (.A(n141[15]), .B(oled_dcn_N_888), .Z(n167[15])) /* synthesis lut_function=(!((B)+!A)) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(88[19:29])
    defparam i13720_2_lut.init = 16'h2222;
    LUT4 mux_414_Mux_27_i15_3_lut_3_lut_4_lut_4_lut (.A(num2[0]), .B(n25753), 
         .C(n25635), .D(n25676), .Z(n23507)) /* synthesis lut_function=(!(A (B (C))+!A (C+!(D)))) */ ;
    defparam mux_414_Mux_27_i15_3_lut_3_lut_4_lut_4_lut.init = 16'h2f2a;
    LUT4 i13719_2_lut (.A(n141[14]), .B(oled_dcn_N_888), .Z(n167[14])) /* synthesis lut_function=(!((B)+!A)) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(88[19:29])
    defparam i13719_2_lut.init = 16'h2222;
    LUT4 i13651_2_lut_3_lut_3_lut_3_lut_4_lut (.A(num2[0]), .B(n25753), 
         .C(n25635), .D(n25676), .Z(n30)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (B+(C+!(D))))) */ ;
    defparam i13651_2_lut_3_lut_3_lut_3_lut_4_lut.init = 16'h0900;
    LUT4 state_0__bdd_4_lut_22149_rep_324 (.A(state[0]), .B(n11_adj_5073), 
         .C(n25684), .D(n25761), .Z(clk_c_enable_1446)) /* synthesis lut_function=(!(A (B (C+!(D)))+!A (B+!(C+!(D))))) */ ;
    defparam state_0__bdd_4_lut_22149_rep_324.init = 16'h3a33;
    LUT4 i13718_2_lut (.A(n141[13]), .B(oled_dcn_N_888), .Z(n167[13])) /* synthesis lut_function=(!((B)+!A)) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(88[19:29])
    defparam i13718_2_lut.init = 16'h2222;
    LUT4 i20778_2_lut_rep_278_3_lut_3_lut_4_lut (.A(num2[0]), .B(n25753), 
         .C(n25676), .D(n25635), .Z(n25560)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (((D)+!C)+!B))) */ ;
    defparam i20778_2_lut_rep_278_3_lut_3_lut_4_lut.init = 16'h0060;
    LUT4 i9227_2_lut_4_lut (.A(state[0]), .B(n11_adj_5073), .C(n25684), 
         .D(n25761), .Z(n12042)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i9227_2_lut_4_lut.init = 16'h0800;
    LUT4 i13717_2_lut (.A(n141[12]), .B(oled_dcn_N_888), .Z(n167[12])) /* synthesis lut_function=(!((B)+!A)) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(88[19:29])
    defparam i13717_2_lut.init = 16'h2222;
    LUT4 state_0__bdd_4_lut_then_4_lut (.A(cnt_scan[2]), .B(cnt_scan[1]), 
         .C(cnt_scan[0]), .D(cnt_scan[3]), .Z(n25788)) /* synthesis lut_function=(A (D)+!A (B (C (D))+!B !((D)+!C))) */ ;
    defparam state_0__bdd_4_lut_then_4_lut.init = 16'hea10;
    LUT4 i13344_2_lut (.A(n141[0]), .B(oled_dcn_N_888), .Z(n167[0])) /* synthesis lut_function=(!((B)+!A)) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(88[19:29])
    defparam i13344_2_lut.init = 16'h2222;
    LUT4 cnt_main_4__bdd_4_lut_22294 (.A(cnt_main[0]), .B(cnt_main[3]), 
         .C(cnt_main[2]), .D(cnt_main[1]), .Z(n24914)) /* synthesis lut_function=(A (B (C))+!A !(B+(C+(D)))) */ ;
    defparam cnt_main_4__bdd_4_lut_22294.init = 16'h8081;
    LUT4 mux_131_Mux_1_i5_3_lut (.A(y_pl[1]), .B(y_ph[1]), .C(cnt_scan[0]), 
         .Z(n5_adj_5048)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(111[7] 142[14])
    defparam mux_131_Mux_1_i5_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_89 (.A(state[2]), .B(n25620), .C(n19), .D(n16_adj_5074), 
         .Z(n6_adj_5075)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_89.init = 16'haaa8;
    LUT4 i13579_2_lut (.A(n25036), .B(cnt_scan[0]), .Z(n6550)) /* synthesis lut_function=(A (B)) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(111[7] 142[14])
    defparam i13579_2_lut.init = 16'h8888;
    LUT4 i13716_2_lut (.A(n141[11]), .B(oled_dcn_N_888), .Z(n167[11])) /* synthesis lut_function=(!((B)+!A)) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(88[19:29])
    defparam i13716_2_lut.init = 16'h2222;
    FD1P3AY y_ph_i0_i1 (.D(n5820[1]), .SP(clk_c_enable_690), .CK(clk_c), 
            .Q(y_ph[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam y_ph_i0_i1.GSR = "ENABLED";
    LUT4 i13715_2_lut (.A(n141[10]), .B(oled_dcn_N_888), .Z(n167[10])) /* synthesis lut_function=(!((B)+!A)) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(88[19:29])
    defparam i13715_2_lut.init = 16'h2222;
    LUT4 i13580_4_lut (.A(cnt_init[0]), .B(n23229), .C(n25581), .D(n25637), 
         .Z(n3871[0])) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i13580_4_lut.init = 16'h0004;
    FD1S3AX x_pl_i3 (.D(x_pl_7__N_529[3]), .CK(clk_c), .Q(x_pl[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam x_pl_i3.GSR = "ENABLED";
    FD1S3AX x_pl_i4 (.D(x_pl_7__N_529[4]), .CK(clk_c), .Q(x_pl[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam x_pl_i4.GSR = "ENABLED";
    FD1S3AX x_pl_i5 (.D(x_pl_7__N_529[5]), .CK(clk_c), .Q(x_pl[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam x_pl_i5.GSR = "ENABLED";
    FD1S3AX x_pl_i6 (.D(x_pl_7__N_529[6]), .CK(clk_c), .Q(x_pl[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam x_pl_i6.GSR = "ENABLED";
    FD1P3AX num1_i0_i3 (.D(n3624[3]), .SP(clk_c_enable_1432), .CK(clk_c), 
            .Q(num1[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam num1_i0_i3.GSR = "ENABLED";
    FD1P3AX num1_i0_i5 (.D(n3624[5]), .SP(clk_c_enable_694), .CK(clk_c), 
            .Q(num1[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam num1_i0_i5.GSR = "ENABLED";
    FD1P3AX num1_i0_i6 (.D(n3624[6]), .SP(clk_c_enable_694), .CK(clk_c), 
            .Q(num1[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam num1_i0_i6.GSR = "ENABLED";
    FD1P3AX num1_i0_i7 (.D(n3624[7]), .SP(clk_c_enable_694), .CK(clk_c), 
            .Q(num1[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam num1_i0_i7.GSR = "ENABLED";
    FD1P3AX num2_i0_i1 (.D(n3536[1]), .SP(clk_c_enable_1431), .CK(clk_c), 
            .Q(num2[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam num2_i0_i1.GSR = "ENABLED";
    FD1P3AX char_reg_i0_i1 (.D(n3492[1]), .SP(clk_c_enable_702), .CK(clk_c), 
            .Q(char_reg[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam char_reg_i0_i1.GSR = "ENABLED";
    FD1P3AX char_reg_i0_i2 (.D(n3492[2]), .SP(clk_c_enable_702), .CK(clk_c), 
            .Q(char_reg[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam char_reg_i0_i2.GSR = "ENABLED";
    FD1P3AX char_reg_i0_i3 (.D(n3492[3]), .SP(clk_c_enable_702), .CK(clk_c), 
            .Q(char_reg[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam char_reg_i0_i3.GSR = "ENABLED";
    FD1P3AX char_reg_i0_i4 (.D(n3492[4]), .SP(clk_c_enable_702), .CK(clk_c), 
            .Q(char_reg[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam char_reg_i0_i4.GSR = "ENABLED";
    FD1P3AX char_reg_i0_i5 (.D(n3492[5]), .SP(clk_c_enable_702), .CK(clk_c), 
            .Q(char_reg[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam char_reg_i0_i5.GSR = "ENABLED";
    FD1P3AX char_reg_i0_i6 (.D(n25040), .SP(clk_c_enable_702), .CK(clk_c), 
            .Q(char_reg[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam char_reg_i0_i6.GSR = "ENABLED";
    FD1P3AX char_reg_i0_i7 (.D(n25191), .SP(clk_c_enable_702), .CK(clk_c), 
            .Q(char_reg[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam char_reg_i0_i7.GSR = "ENABLED";
    FD1S3AX char_i1 (.D(char_7__N_553[1]), .CK(clk_c), .Q(char[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam char_i1.GSR = "ENABLED";
    FD1S3AX char_i2 (.D(char_7__N_553[2]), .CK(clk_c), .Q(char[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam char_i2.GSR = "ENABLED";
    FD1S3AX char_i3 (.D(char_7__N_553[3]), .CK(clk_c), .Q(char[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam char_i3.GSR = "ENABLED";
    FD1S3AX char_i4 (.D(char_7__N_553[4]), .CK(clk_c), .Q(char[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam char_i4.GSR = "ENABLED";
    FD1S3AX char_i5 (.D(char_7__N_553[5]), .CK(clk_c), .Q(char[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam char_i5.GSR = "ENABLED";
    FD1S3AX char_i6 (.D(char_7__N_553[6]), .CK(clk_c), .Q(char[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam char_i6.GSR = "ENABLED";
    FD1S3AX num1_delay_i1 (.D(num1_delay_15__N_605[1]), .CK(clk_c), .Q(num1_delay[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam num1_delay_i1.GSR = "ENABLED";
    FD1S3AY num1_delay_i2 (.D(num1_delay_15__N_605[2]), .CK(clk_c), .Q(num1_delay[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam num1_delay_i2.GSR = "ENABLED";
    FD1S3AX num1_delay_i3 (.D(num1_delay_15__N_605[3]), .CK(clk_c), .Q(num1_delay[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam num1_delay_i3.GSR = "ENABLED";
    FD1S3AX num1_delay_i4 (.D(num1_delay_15__N_605[4]), .CK(clk_c), .Q(num1_delay[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam num1_delay_i4.GSR = "ENABLED";
    FD1S3AX num1_delay_i5 (.D(num1_delay_15__N_605[5]), .CK(clk_c), .Q(num1_delay[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam num1_delay_i5.GSR = "ENABLED";
    FD1S3AX num1_delay_i6 (.D(num1_delay_15__N_605[6]), .CK(clk_c), .Q(num1_delay[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam num1_delay_i6.GSR = "ENABLED";
    FD1S3AX num1_delay_i7 (.D(num1_delay_15__N_605[7]), .CK(clk_c), .Q(num1_delay[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam num1_delay_i7.GSR = "ENABLED";
    FD1S3AX num1_delay_i8 (.D(num1_delay_15__N_605[8]), .CK(clk_c), .Q(num1_delay[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam num1_delay_i8.GSR = "ENABLED";
    FD1S3AX num1_delay_i9 (.D(num1_delay_15__N_605[9]), .CK(clk_c), .Q(num1_delay[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam num1_delay_i9.GSR = "ENABLED";
    FD1S3AX num1_delay_i10 (.D(num1_delay_15__N_605[10]), .CK(clk_c), .Q(num1_delay[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam num1_delay_i10.GSR = "ENABLED";
    FD1S3AX num1_delay_i11 (.D(num1_delay_15__N_605[11]), .CK(clk_c), .Q(num1_delay[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam num1_delay_i11.GSR = "ENABLED";
    FD1S3AX num1_delay_i12 (.D(num1_delay_15__N_605[12]), .CK(clk_c), .Q(num1_delay[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam num1_delay_i12.GSR = "ENABLED";
    FD1S3AX num1_delay_i13 (.D(num1_delay_15__N_605[13]), .CK(clk_c), .Q(num1_delay[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam num1_delay_i13.GSR = "ENABLED";
    FD1S3AX num1_delay_i14 (.D(num1_delay_15__N_605[14]), .CK(clk_c), .Q(num1_delay[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam num1_delay_i14.GSR = "ENABLED";
    FD1S3AX num1_delay_i15 (.D(num1_delay_15__N_605[15]), .CK(clk_c), .Q(num1_delay[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam num1_delay_i15.GSR = "ENABLED";
    FD1S3AX state_back_i1 (.D(state_back_5__N_659[1]), .CK(clk_c), .Q(state_back[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam state_back_i1.GSR = "ENABLED";
    FD1S3AX state_back_i2 (.D(state_back_5__N_659[2]), .CK(clk_c), .Q(state_back[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam state_back_i2.GSR = "ENABLED";
    FD1S3AX state_back_i3 (.D(state_back_5__N_659[3]), .CK(clk_c), .Q(state_back[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam state_back_i3.GSR = "ENABLED";
    FD1S3AX state_back_i4 (.D(state_back_5__N_659[4]), .CK(clk_c), .Q(state_back[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam state_back_i4.GSR = "ENABLED";
    FD1S3AX state_back_i5 (.D(state_back_5__N_659[5]), .CK(clk_c), .Q(state_back[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam state_back_i5.GSR = "ENABLED";
    FD1S3AY x_ph_i1 (.D(x_ph_7__N_519[1]), .CK(clk_c), .Q(x_ph[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam x_ph_i1.GSR = "ENABLED";
    FD1S3AY x_ph_i2 (.D(x_ph_7__N_519[2]), .CK(clk_c), .Q(x_ph[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam x_ph_i2.GSR = "ENABLED";
    FD1S3AY x_ph_i3 (.D(x_ph_7__N_519[3]), .CK(clk_c), .Q(x_ph[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam x_ph_i3.GSR = "ENABLED";
    FD1S3AY x_ph_i4 (.D(x_ph_7__N_519[4]), .CK(clk_c), .Q(x_ph[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam x_ph_i4.GSR = "ENABLED";
    FD1S3AY x_ph_i5 (.D(x_ph_7__N_519[5]), .CK(clk_c), .Q(x_ph[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam x_ph_i5.GSR = "ENABLED";
    FD1S3AY x_ph_i6 (.D(x_ph_7__N_519[6]), .CK(clk_c), .Q(x_ph[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam x_ph_i6.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_4_lut_adj_90 (.A(cnt_main[1]), .B(n25743), .C(char[6]), 
         .D(cnt_main[4]), .Z(n43_adj_5076)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_90.init = 16'hf080;
    LUT4 i13714_2_lut (.A(n141[9]), .B(oled_dcn_N_888), .Z(n167[9])) /* synthesis lut_function=(!((B)+!A)) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(88[19:29])
    defparam i13714_2_lut.init = 16'h2222;
    LUT4 i1_2_lut_3_lut_4_lut_adj_91 (.A(cnt_main[1]), .B(n25743), .C(x_pl[5]), 
         .D(cnt_main[4]), .Z(n27_adj_5077)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_91.init = 16'hf080;
    LUT4 i13713_2_lut (.A(n141[8]), .B(oled_dcn_N_888), .Z(n167[8])) /* synthesis lut_function=(!((B)+!A)) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(88[19:29])
    defparam i13713_2_lut.init = 16'h2222;
    LUT4 i3_4_lut_adj_92 (.A(num2[0]), .B(n25686), .C(n6178), .D(n16320), 
         .Z(n20729)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(111[7] 142[14])
    defparam i3_4_lut_adj_92.init = 16'h0020;
    PFUMX i21667 (.BLUT(n24714), .ALUT(n24713), .C0(cnt_main[3]), .Z(n24715));
    LUT4 i1_2_lut_4_lut (.A(n25745), .B(char[4]), .C(char[3]), .D(char[5]), 
         .Z(n23153)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(129[56:62])
    defparam i1_2_lut_4_lut.init = 16'h8000;
    LUT4 i13712_2_lut (.A(n141[7]), .B(oled_dcn_N_888), .Z(n167[7])) /* synthesis lut_function=(!((B)+!A)) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(88[19:29])
    defparam i13712_2_lut.init = 16'h2222;
    LUT4 i1_3_lut_4_lut (.A(n25750), .B(n25749), .C(n9), .D(x_ph[5]), 
         .Z(n4_adj_5078)) /* synthesis lut_function=(!(A (C (D))+!A ((C (D))+!B))) */ ;
    defparam i1_3_lut_4_lut.init = 16'h0eee;
    LUT4 i13711_2_lut (.A(n141[6]), .B(oled_dcn_N_888), .Z(n167[6])) /* synthesis lut_function=(!((B)+!A)) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(88[19:29])
    defparam i13711_2_lut.init = 16'h2222;
    LUT4 i24_3_lut_4_lut (.A(state[0]), .B(n25646), .C(state[1]), .D(n12_adj_5079), 
         .Z(n22465)) /* synthesis lut_function=(A (B (D)+!B ((D)+!C))+!A (B (D)+!B !(C+!(D)))) */ ;
    defparam i24_3_lut_4_lut.init = 16'hef02;
    LUT4 i1_2_lut_3_lut_4_lut_adj_93 (.A(cnt_main[4]), .B(n25744), .C(state[1]), 
         .D(n25750), .Z(n5_adj_5080)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_93.init = 16'h0010;
    LUT4 i13710_2_lut (.A(n141[5]), .B(oled_dcn_N_888), .Z(n167[5])) /* synthesis lut_function=(!((B)+!A)) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(88[19:29])
    defparam i13710_2_lut.init = 16'h2222;
    LUT4 i2_3_lut_adj_94 (.A(state[1]), .B(state[2]), .C(state[0]), .Z(n8)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(77[5:9])
    defparam i2_3_lut_adj_94.init = 16'hfbfb;
    LUT4 i13709_2_lut (.A(n141[4]), .B(oled_dcn_N_888), .Z(n167[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(88[19:29])
    defparam i13709_2_lut.init = 16'h2222;
    LUT4 i13708_2_lut (.A(n141[3]), .B(oled_dcn_N_888), .Z(n167[3])) /* synthesis lut_function=(!((B)+!A)) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(88[19:29])
    defparam i13708_2_lut.init = 16'h2222;
    LUT4 i21284_3_lut (.A(n26455), .B(n23350), .C(cnt_scan[3]), .Z(n23898)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21284_3_lut.init = 16'hcaca;
    LUT4 i13707_2_lut (.A(n141[2]), .B(oled_dcn_N_888), .Z(n167[2])) /* synthesis lut_function=(!((B)+!A)) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(88[19:29])
    defparam i13707_2_lut.init = 16'h2222;
    LUT4 i1_2_lut_3_lut_4_lut_adj_95 (.A(n25691), .B(n25649), .C(n25636), 
         .D(n25692), .Z(n4_adj_5081)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A ((D)+!C))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_95.init = 16'h00d0;
    LUT4 i20895_4_lut (.A(num2[0]), .B(n23694), .C(n25074), .D(cnt_scan[0]), 
         .Z(n23769)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i20895_4_lut.init = 16'ha088;
    LUT4 i21055_3_lut (.A(n23930), .B(n23931), .C(cnt_scan[2]), .Z(n23932)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21055_3_lut.init = 16'hcaca;
    LUT4 i21289_3_lut (.A(n23932), .B(n23769), .C(cnt_scan[3]), .Z(n23907)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21289_3_lut.init = 16'hcaca;
    LUT4 i13706_2_lut (.A(n141[1]), .B(oled_dcn_N_888), .Z(n167[1])) /* synthesis lut_function=(!((B)+!A)) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(88[19:29])
    defparam i13706_2_lut.init = 16'h2222;
    LUT4 state_0__bdd_4_lut_else_4_lut (.A(cnt_scan[2]), .B(cnt_scan[1]), 
         .C(cnt_scan[0]), .D(cnt_scan[3]), .Z(n25787)) /* synthesis lut_function=(A (D)+!A (B (C (D)))) */ ;
    defparam state_0__bdd_4_lut_else_4_lut.init = 16'hea00;
    LUT4 i21020_4_lut (.A(n6), .B(n23920), .C(cnt_scan[3]), .D(cnt_scan[2]), 
         .Z(n23897)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam i21020_4_lut.init = 16'hcac0;
    LUT4 mux_131_Mux_2_i22_4_lut (.A(n18_adj_5082), .B(n25316), .C(cnt_scan[2]), 
         .D(cnt_scan[0]), .Z(n22)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(111[7] 142[14])
    defparam mux_131_Mux_2_i22_4_lut.init = 16'hca0a;
    LUT4 i21295_3_lut (.A(n22), .B(n23348), .C(cnt_scan[3]), .Z(n23895)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21295_3_lut.init = 16'hcaca;
    PFUMX i21665 (.BLUT(n24711), .ALUT(n24710), .C0(cnt_scan[2]), .Z(n24712));
    LUT4 i21557_2_lut_3_lut_3_lut (.A(n25601), .B(cnt_scan[0]), .C(n25635), 
         .Z(n23867)) /* synthesis lut_function=(((C)+!B)+!A) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(111[7] 142[14])
    defparam i21557_2_lut_3_lut_3_lut.init = 16'hf7f7;
    LUT4 i21037_3_lut (.A(n25216), .B(n23913), .C(cnt_scan[2]), .Z(n23914)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21037_3_lut.init = 16'hcaca;
    FD1P3IX cnt_scan_i0_i4 (.D(cnt_scan_4__N_682[4]), .SP(clk_c_enable_1446), 
            .CD(n12042), .CK(clk_c), .Q(cnt_scan[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam cnt_scan_i0_i4.GSR = "ENABLED";
    FD1P3IX cnt_scan_i0_i3 (.D(cnt_scan_4__N_682[3]), .SP(clk_c_enable_1446), 
            .CD(n12042), .CK(clk_c), .Q(cnt_scan[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam cnt_scan_i0_i3.GSR = "ENABLED";
    FD1P3IX cnt_scan_i0_i1 (.D(cnt_scan_4__N_682[1]), .SP(clk_c_enable_1446), 
            .CD(n12042), .CK(clk_c), .Q(cnt_scan[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam cnt_scan_i0_i1.GSR = "ENABLED";
    FD1P3IX cnt_main_1988__i4 (.D(n25771), .SP(clk_c_enable_1352), .CD(n12039), 
            .CK(clk_c), .Q(cnt_main[4]));   // g:/fpga/mxo2/system/project/oled12832.v(53[12:40])
    defparam cnt_main_1988__i4.GSR = "ENABLED";
    LUT4 i21297_3_lut (.A(n23914), .B(n26778), .C(cnt_scan[3]), .Z(n23892)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21297_3_lut.init = 16'hcaca;
    LUT4 i20668_2_lut_rep_342_4_lut (.A(num2[2]), .B(char[2]), .C(n25752), 
         .D(num2[0]), .Z(n25624)) /* synthesis lut_function=(A (B (C+(D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C+(D)))) */ ;
    defparam i20668_2_lut_rep_342_4_lut.init = 16'hff96;
    LUT4 n25425_bdd_4_lut_then_4_lut (.A(cnt_main[3]), .B(cnt_main[4]), 
         .C(cnt_main[0]), .D(cnt_main[1]), .Z(n25791)) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A (B+(D)))) */ ;
    defparam n25425_bdd_4_lut_then_4_lut.init = 16'h0211;
    LUT4 n25425_bdd_4_lut_else_4_lut (.A(cnt_main[3]), .B(cnt_main[4]), 
         .C(cnt_main[0]), .D(cnt_main[1]), .Z(n25790)) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam n25425_bdd_4_lut_else_4_lut.init = 16'h1110;
    LUT4 i1_2_lut_adj_96 (.A(state[2]), .B(state[0]), .Z(n23590)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_96.init = 16'h8888;
    LUT4 i20886_2_lut (.A(cnt_init[2]), .B(cnt_init[1]), .Z(n23755)) /* synthesis lut_function=(A (B)) */ ;
    defparam i20886_2_lut.init = 16'h8888;
    LUT4 i21029_3_lut (.A(n24712), .B(n23941), .C(cnt_scan[3]), .Z(n23906)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21029_3_lut.init = 16'hcaca;
    LUT4 i2_4_lut_adj_97 (.A(n4_adj_5083), .B(n4_adj_5081), .C(state[0]), 
         .D(n25608), .Z(clk_c_enable_1421)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i2_4_lut_adj_97.init = 16'hc088;
    PFUMX i21656 (.BLUT(n24696), .ALUT(n24695), .C0(cnt_main[0]), .Z(n24697));
    LUT4 i2_3_lut_adj_98 (.A(cnt_write[4]), .B(state[4]), .C(cnt_write[0]), 
         .Z(n4_adj_5083)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i2_3_lut_adj_98.init = 16'h4040;
    PFUMX i21922 (.BLUT(n25553), .ALUT(n25189), .C0(state[3]), .Z(n25191));
    LUT4 i2_3_lut_adj_99 (.A(n25608), .B(state[4]), .C(n23881), .Z(n20727)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(27[43:52])
    defparam i2_3_lut_adj_99.init = 16'h4040;
    LUT4 i13530_2_lut (.A(num2[0]), .B(n25121), .Z(n23_adj_5084)) /* synthesis lut_function=(A (B)) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(111[7] 142[14])
    defparam i13530_2_lut.init = 16'h8888;
    LUT4 i21050_4_lut (.A(n16_adj_5085), .B(n23716), .C(cnt_scan[1]), 
         .D(n23422), .Z(n23927)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam i21050_4_lut.init = 16'h0aca;
    LUT4 i21052_3_lut (.A(n23927), .B(n23928), .C(cnt_scan[2]), .Z(n23929)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21052_3_lut.init = 16'hcaca;
    LUT4 i21299_3_lut (.A(n23929), .B(n23_adj_5084), .C(cnt_scan[3]), 
         .Z(n23904)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21299_3_lut.init = 16'hcaca;
    LUT4 i21023_3_lut (.A(n7), .B(n23923), .C(cnt_scan[3]), .Z(n23900)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21023_3_lut.init = 16'hcaca;
    LUT4 i4306_3_lut_4_lut_4_lut (.A(n25601), .B(n24966), .C(n25594), 
         .D(n25667), .Z(n7109)) /* synthesis lut_function=(A (B)+!A (C (D))) */ ;
    defparam i4306_3_lut_4_lut_4_lut.init = 16'hd888;
    FD1P3IX cnt_main_1988__i3 (.D(n25872), .SP(clk_c_enable_1352), .CD(n12039), 
            .CK(clk_c), .Q(cnt_main[3]));   // g:/fpga/mxo2/system/project/oled12832.v(53[12:40])
    defparam cnt_main_1988__i3.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_100 (.A(n21029), .B(n25751), .C(n6_adj_5086), .D(cnt[3]), 
         .Z(oled_dcn_N_888)) /* synthesis lut_function=(A+!(B+!(C (D)))) */ ;
    defparam i1_4_lut_adj_100.init = 16'hbaaa;
    LUT4 i21017_4_lut (.A(cnt_scan[2]), .B(n23917), .C(cnt_scan[3]), .D(n4_adj_5087), 
         .Z(n23894)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam i21017_4_lut.init = 16'hcac0;
    LUT4 n24965_bdd_3_lut_4_lut (.A(n25753), .B(num2[0]), .C(cnt_scan[0]), 
         .D(n24964), .Z(n24966)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B (C (D))+!B ((D)+!C))) */ ;
    defparam n24965_bdd_3_lut_4_lut.init = 16'hf909;
    LUT4 i21014_3_lut (.A(n24683), .B(n23911), .C(cnt_scan[3]), .Z(n23891)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21014_3_lut.init = 16'hcaca;
    LUT4 i17716_3_lut (.A(char[3]), .B(num2[3]), .C(n6_adj_5088), .Z(n8_adj_5054)) /* synthesis lut_function=(A ((C)+!B)+!A !(B+!(C))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(139[77:83])
    defparam i17716_3_lut.init = 16'hb2b2;
    LUT4 i1_3_lut (.A(n20788), .B(n83), .C(x_ph[0]), .Z(x_ph_7__N_519[0])) /* synthesis lut_function=(!(A (B)+!A !((C)+!B))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(29[13:18])
    defparam i1_3_lut.init = 16'h7373;
    LUT4 i21418_3_lut_rep_299_4_lut (.A(n25756), .B(n25755), .C(cnt_init[0]), 
         .D(oled_dcn_N_888), .Z(n25581)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(92[8:12])
    defparam i21418_3_lut_rep_299_4_lut.init = 16'h0001;
    LUT4 i4_4_lut (.A(state[0]), .B(n89), .C(n58), .D(n6_adj_5089), 
         .Z(n20788)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i4_4_lut.init = 16'h4000;
    LUT4 i21026_3_lut (.A(n7_adj_5060), .B(n23926), .C(cnt_scan[3]), .Z(n23903)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21026_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_4_lut (.A(n25756), .B(n25755), .C(n23755), .D(cnt_init[0]), 
         .Z(n23229)) /* synthesis lut_function=(!(A+(B (C)+!B (C+(D))))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(92[8:12])
    defparam i1_4_lut_4_lut.init = 16'h0405;
    LUT4 i10_4_lut (.A(cnt_c[5]), .B(n20), .C(n16_adj_5090), .D(cnt_c[10]), 
         .Z(n21029)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i10_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_adj_101 (.A(state[1]), .B(cnt_main[4]), .Z(n6_adj_5089)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut_adj_101.init = 16'h2222;
    LUT4 i4271_3_lut_rep_304_4_lut (.A(cnt_scan[3]), .B(n25660), .C(cnt_scan[4]), 
         .D(n8418), .Z(n25586)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A (C (D)))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(111[7] 142[14])
    defparam i4271_3_lut_rep_304_4_lut.init = 16'h0dfd;
    LUT4 i1_4_lut_adj_102 (.A(state[0]), .B(x_pl[3]), .C(n16_adj_5091), 
         .D(n19_adj_5092), .Z(x_pl_7__N_529[3])) /* synthesis lut_function=(A (B (D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_102.init = 16'hdc50;
    PFUMX i21919 (.BLUT(n25186), .ALUT(n20729), .C0(cnt_scan[3]), .Z(n25187));
    LUT4 i33_4_lut (.A(x_pl[3]), .B(x_pl_7__N_700[3]), .C(state[1]), .D(n25646), 
         .Z(n16_adj_5091)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam i33_4_lut.init = 16'h0aca;
    LUT4 i2_2_lut_adj_103 (.A(cnt[4]), .B(cnt[2]), .Z(n6_adj_5086)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2_2_lut_adj_103.init = 16'h8888;
    LUT4 i1_4_lut_adj_104 (.A(n19_adj_5092), .B(state[1]), .C(state[0]), 
         .D(n89), .Z(n83)) /* synthesis lut_function=(A+!(B (C+!(D))+!B (C))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(29[13:18])
    defparam i1_4_lut_adj_104.init = 16'hafab;
    LUT4 i2_4_lut_adj_105 (.A(n25578), .B(n15856), .C(x_pl[3]), .D(n9), 
         .Z(x_pl_7__N_700[3])) /* synthesis lut_function=(((C (D))+!B)+!A) */ ;
    defparam i2_4_lut_adj_105.init = 16'hf777;
    LUT4 i9_4_lut (.A(cnt_c[9]), .B(n18_adj_5093), .C(cnt_c[8]), .D(cnt_c[6]), 
         .Z(n20)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i9_4_lut.init = 16'hfffe;
    LUT4 i2_4_lut_adj_106 (.A(n25115), .B(n4_adj_5094), .C(state[0]), 
         .D(n25608), .Z(clk_c_enable_1423)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i2_4_lut_adj_106.init = 16'hc088;
    LUT4 i2_4_lut_adj_107 (.A(n25682), .B(state[4]), .C(cnt_write[4]), 
         .D(cnt_write[0]), .Z(n12_adj_5079)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (((D)+!C)+!B))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(41[4] 175[11])
    defparam i2_4_lut_adj_107.init = 16'h0048;
    LUT4 i5_2_lut (.A(cnt_c[11]), .B(cnt_c[13]), .Z(n16_adj_5090)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i5_2_lut.init = 16'heeee;
    LUT4 i1_4_lut_adj_108 (.A(state[1]), .B(n20715), .C(n23718), .D(state[5]), 
         .Z(n3264)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B+!(C+!(D)))) */ ;
    defparam i1_4_lut_adj_108.init = 16'hcdce;
    LUT4 i7_4_lut_adj_109 (.A(cnt_c[7]), .B(cnt_c[14]), .C(cnt_c[12]), 
         .D(cnt_c[15]), .Z(n18_adj_5093)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut_adj_109.init = 16'hfffe;
    LUT4 i21574_3_lut_3_lut_4_lut (.A(state[2]), .B(n25684), .C(n10049), 
         .D(n25683), .Z(clk_c_enable_1352)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i21574_3_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i2_3_lut_rep_305_4_lut (.A(state[2]), .B(n25684), .C(state[1]), 
         .D(state[0]), .Z(n25587)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;
    defparam i2_3_lut_rep_305_4_lut.init = 16'hffef;
    LUT4 i1_2_lut_adj_110 (.A(cnt_scan[0]), .B(num2[0]), .Z(n23347)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_110.init = 16'h8888;
    PFUMX i22153 (.BLUT(n25769), .ALUT(n25770), .C0(cnt_main[3]), .Z(n25771));
    LUT4 i1_4_lut_adj_111 (.A(state[0]), .B(x_pl[4]), .C(n16_adj_5095), 
         .D(n19_adj_5092), .Z(x_pl_7__N_529[4])) /* synthesis lut_function=(A (B (D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_111.init = 16'hdc50;
    LUT4 i33_4_lut_adj_112 (.A(x_pl[4]), .B(x_pl_7__N_700[4]), .C(state[1]), 
         .D(n25646), .Z(n16_adj_5095)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam i33_4_lut_adj_112.init = 16'h0aca;
    LUT4 i1_4_lut_adj_113 (.A(n25578), .B(x_pl[4]), .C(n4_adj_5096), .D(n25631), 
         .Z(x_pl_7__N_700[4])) /* synthesis lut_function=((B (C+(D))+!B (C))+!A) */ ;
    defparam i1_4_lut_adj_113.init = 16'hfdf5;
    LUT4 i21053_4_lut (.A(n16_adj_5085), .B(num2[0]), .C(cnt_scan[1]), 
         .D(n8723), .Z(n23930)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (B+((D)+!C)))) */ ;
    defparam i21053_4_lut.init = 16'h0a3a;
    LUT4 i1_4_lut_adj_114 (.A(state[0]), .B(x_pl[5]), .C(n16_adj_5097), 
         .D(n19_adj_5092), .Z(x_pl_7__N_529[5])) /* synthesis lut_function=(A (B (D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_114.init = 16'hdc50;
    LUT4 i33_4_lut_adj_115 (.A(x_pl[5]), .B(x_pl_7__N_700[5]), .C(state[1]), 
         .D(n25646), .Z(n16_adj_5097)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam i33_4_lut_adj_115.init = 16'h0aca;
    LUT4 i1_4_lut_adj_116 (.A(n15856), .B(n5_adj_5098), .C(n25674), .D(n27_adj_5077), 
         .Z(x_pl_7__N_700[5])) /* synthesis lut_function=((B+((D)+!C))+!A) */ ;
    defparam i1_4_lut_adj_116.init = 16'hffdf;
    LUT4 i1_4_lut_adj_117 (.A(cnt_main[0]), .B(n20_adj_5099), .C(n25073), 
         .D(n15942), .Z(n5_adj_5098)) /* synthesis lut_function=(!(A ((D)+!B)+!A !(B (C+!(D))+!B (C)))) */ ;
    defparam i1_4_lut_adj_117.init = 16'h50dc;
    LUT4 i1_4_lut_4_lut_adj_118 (.A(n25601), .B(n25564), .C(n23347), .D(n25575), 
         .Z(n23349)) /* synthesis lut_function=(A (C (D))+!A !(B+!(C))) */ ;
    defparam i1_4_lut_4_lut_adj_118.init = 16'hb010;
    LUT4 i13167_2_lut (.A(cnt_main[4]), .B(cnt_main[3]), .Z(n15942)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i13167_2_lut.init = 16'heeee;
    FD1P3IX cnt_main_1988__i2 (.D(n23589), .SP(clk_c_enable_1352), .CD(n12039), 
            .CK(clk_c), .Q(cnt_main[2]));   // g:/fpga/mxo2/system/project/oled12832.v(53[12:40])
    defparam cnt_main_1988__i2.GSR = "ENABLED";
    LUT4 i1_4_lut_4_lut_adj_119 (.A(n25601), .B(n23803), .C(n23347), .D(n25575), 
         .Z(n23350)) /* synthesis lut_function=(A (C (D))+!A (B (C))) */ ;
    defparam i1_4_lut_4_lut_adj_119.init = 16'he040;
    LUT4 i1_4_lut_adj_120 (.A(state[0]), .B(n19_adj_5092), .C(n17773), 
         .D(x_pl[6]), .Z(x_pl_7__N_529[6])) /* synthesis lut_function=(A (B (D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_120.init = 16'hdc50;
    LUT4 i1_3_lut_adj_121 (.A(cnt_main[2]), .B(cnt_main[0]), .C(time_data[3]), 
         .Z(n86)) /* synthesis lut_function=(A (B+!(C))) */ ;
    defparam i1_3_lut_adj_121.init = 16'h8a8a;
    LUT4 i2737_3_lut_4_lut (.A(cnt_write[2]), .B(n25758), .C(cnt_write[3]), 
         .D(cnt_write[4]), .Z(n2535[4])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(146[25:41])
    defparam i2737_3_lut_4_lut.init = 16'h7f80;
    LUT4 i15050_4_lut (.A(x_pl[6]), .B(n23159), .C(state[1]), .D(n25646), 
         .Z(n17773)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (B+((D)+!C)))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(29[13:18])
    defparam i15050_4_lut.init = 16'h0a3a;
    LUT4 i1_4_lut_adj_122 (.A(n60), .B(n23157), .C(x_pl[6]), .D(n62_adj_5100), 
         .Z(n23159)) /* synthesis lut_function=(A (B)+!A !((C+!(D))+!B)) */ ;
    defparam i1_4_lut_adj_122.init = 16'h8c88;
    LUT4 i2357_2_lut_rep_356_4_lut (.A(cnt_write[1]), .B(n25694), .C(cnt_write[4]), 
         .D(cnt_write[0]), .Z(n25638)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(147[7] 167[14])
    defparam i2357_2_lut_rep_356_4_lut.init = 16'hf0e0;
    LUT4 mux_1293_i4_4_lut (.A(num1_7__N_724[3]), .B(num1_7__N_732[3]), 
         .C(state[3]), .D(state[0]), .Z(n3624[3])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;
    defparam mux_1293_i4_4_lut.init = 16'hc0ca;
    LUT4 i1_4_lut_adj_123 (.A(n29), .B(state[3]), .C(n16391), .D(n25585), 
         .Z(clk_c_enable_694)) /* synthesis lut_function=(!((B ((D)+!C)+!B !(C))+!A)) */ ;
    defparam i1_4_lut_adj_123.init = 16'h20a0;
    LUT4 i20992_2_lut (.A(n1354), .B(n1355), .Z(n23869)) /* synthesis lut_function=(!(A+!(B))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(129[51:75])
    defparam i20992_2_lut.init = 16'h4444;
    LUT4 i21335_4_lut (.A(n16678), .B(n24049), .C(n4432), .D(n25609), 
         .Z(clk_c_enable_1427)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A !(B (C+(D))))) */ ;
    defparam i21335_4_lut.init = 16'h44c0;
    LUT4 i49_4_lut (.A(cnt_scan[4]), .B(n25581), .C(state[2]), .D(n8418), 
         .Z(n16678)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (B+!(C)))) */ ;
    defparam i49_4_lut.init = 16'h3a30;
    LUT4 i21334_4_lut (.A(n25660), .B(n3264), .C(n6_adj_5101), .D(cnt_scan[4]), 
         .Z(n24049)) /* synthesis lut_function=(A (B)+!A (B ((D)+!C))) */ ;
    defparam i21334_4_lut.init = 16'hcc8c;
    LUT4 i2_3_lut_4_lut (.A(state[0]), .B(n25761), .C(n25760), .D(state[3]), 
         .Z(n11_adj_5073)) /* synthesis lut_function=(A+((C+!(D))+!B)) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(169[5:10])
    defparam i2_3_lut_4_lut.init = 16'hfbff;
    LUT4 i13330_2_lut_rep_296_3_lut_4_lut (.A(cnt_main[3]), .B(n25658), 
         .C(n25711), .D(n25718), .Z(n25578)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B !(C))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(59[8:12])
    defparam i13330_2_lut_rep_296_3_lut_4_lut.init = 16'hef0f;
    LUT4 i21426_3_lut_4_lut (.A(state[0]), .B(n25761), .C(n25684), .D(n24139), 
         .Z(clk_c_enable_1359)) /* synthesis lut_function=(!(A (C+!(D))+!A (B+(C+!(D))))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(169[5:10])
    defparam i21426_3_lut_4_lut.init = 16'h0b00;
    LUT4 mux_1262_i2_4_lut (.A(n25657), .B(num2_7__N_748[1]), .C(state[3]), 
         .D(state[0]), .Z(n3536[1])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;
    defparam mux_1262_i2_4_lut.init = 16'hc0ca;
    LUT4 i1_4_lut_adj_124 (.A(n25660), .B(n25593), .C(cnt_scan[4]), .D(cnt_scan[3]), 
         .Z(n23342)) /* synthesis lut_function=(A (B (C+(D)))+!A (B (C))) */ ;
    defparam i1_4_lut_adj_124.init = 16'hc8c0;
    LUT4 mux_1250_i2_4_lut (.A(n25558), .B(char_reg_7__N_772[1]), .C(state[3]), 
         .D(n25539), .Z(n3492[1])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_1250_i2_4_lut.init = 16'hcac0;
    FD1P3IX cnt_main_1988__i1 (.D(n25799), .SP(clk_c_enable_1352), .CD(n12039), 
            .CK(clk_c), .Q(cnt_main[1]));   // g:/fpga/mxo2/system/project/oled12832.v(53[12:40])
    defparam cnt_main_1988__i1.GSR = "ENABLED";
    LUT4 mux_1250_i3_4_lut (.A(n23974), .B(char_reg_7__N_772[2]), .C(state[3]), 
         .D(n25558), .Z(n3492[2])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_1250_i3_4_lut.init = 16'hcac0;
    LUT4 mux_1250_i4_4_lut (.A(n23971), .B(char_reg_7__N_772[3]), .C(state[3]), 
         .D(n25558), .Z(n3492[3])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_1250_i4_4_lut.init = 16'hcac0;
    LUT4 mux_1250_i5_4_lut (.A(n22685), .B(char_reg_7__N_772[4]), .C(state[3]), 
         .D(n25558), .Z(n3492[4])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_1250_i5_4_lut.init = 16'hcac0;
    LUT4 i2665_3_lut_4_lut (.A(cnt_init[2]), .B(n25759), .C(cnt_init[3]), 
         .D(cnt_init[4]), .Z(n1[4])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(79[49:64])
    defparam i2665_3_lut_4_lut.init = 16'h7f80;
    CCU2D add_143_17 (.A0(cnt_delay[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n20504), .S0(n2559[15]));   // g:/fpga/mxo2/system/project/oled12832.v(172[29:45])
    defparam add_143_17.INIT0 = 16'h5aaa;
    defparam add_143_17.INIT1 = 16'h0000;
    defparam add_143_17.INJECT1_0 = "NO";
    defparam add_143_17.INJECT1_1 = "NO";
    CCU2D sub_1361_add_2_17 (.A0(cnt_delay[15]), .B0(num1_delay[15]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n20592), .S1(n2557));
    defparam sub_1361_add_2_17.INIT0 = 16'h5999;
    defparam sub_1361_add_2_17.INIT1 = 16'h0000;
    defparam sub_1361_add_2_17.INJECT1_0 = "NO";
    defparam sub_1361_add_2_17.INJECT1_1 = "NO";
    LUT4 mux_1250_i6_4_lut (.A(n25774), .B(char_reg_7__N_772[5]), .C(state[3]), 
         .D(n25558), .Z(n3492[5])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mux_1250_i6_4_lut.init = 16'hcac0;
    LUT4 i33_4_lut_adj_125 (.A(state[4]), .B(state[0]), .C(n25608), .D(n23223), 
         .Z(n20_adj_5102)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam i33_4_lut_adj_125.init = 16'hcac0;
    LUT4 i2_2_lut_3_lut_3_lut_4_lut (.A(state[3]), .B(n25760), .C(n25761), 
         .D(state[0]), .Z(n12039)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(77[5:9])
    defparam i2_2_lut_3_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i1_3_lut_4_lut_adj_126 (.A(cnt_init[0]), .B(n25677), .C(n25650), 
         .D(num1_delay[7]), .Z(n4_adj_5103)) /* synthesis lut_function=(A ((C (D))+!B)+!A (C (D))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam i1_3_lut_4_lut_adj_126.init = 16'hf222;
    FD1P3IX cnt_init_i0_i1 (.D(n1[1]), .SP(clk_c_enable_1359), .CD(n12024), 
            .CK(clk_c), .Q(cnt_init[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam cnt_init_i0_i1.GSR = "ENABLED";
    CCU2D sub_1361_add_2_15 (.A0(cnt_delay[13]), .B0(num1_delay[13]), .C0(GND_net), 
          .D0(GND_net), .A1(cnt_delay[14]), .B1(num1_delay[14]), .C1(GND_net), 
          .D1(GND_net), .CIN(n20591), .COUT(n20592));
    defparam sub_1361_add_2_15.INIT0 = 16'h5999;
    defparam sub_1361_add_2_15.INIT1 = 16'h5999;
    defparam sub_1361_add_2_15.INJECT1_0 = "NO";
    defparam sub_1361_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_1361_add_2_13 (.A0(cnt_delay[11]), .B0(num1_delay[11]), .C0(GND_net), 
          .D0(GND_net), .A1(cnt_delay[12]), .B1(num1_delay[12]), .C1(GND_net), 
          .D1(GND_net), .CIN(n20590), .COUT(n20591));
    defparam sub_1361_add_2_13.INIT0 = 16'h5999;
    defparam sub_1361_add_2_13.INIT1 = 16'h5999;
    defparam sub_1361_add_2_13.INJECT1_0 = "NO";
    defparam sub_1361_add_2_13.INJECT1_1 = "NO";
    CCU2D add_143_15 (.A0(cnt_delay[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt_delay[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n20503), .COUT(n20504), .S0(n2559[13]), 
          .S1(n2559[14]));   // g:/fpga/mxo2/system/project/oled12832.v(172[29:45])
    defparam add_143_15.INIT0 = 16'h5aaa;
    defparam add_143_15.INIT1 = 16'h5aaa;
    defparam add_143_15.INJECT1_0 = "NO";
    defparam add_143_15.INJECT1_1 = "NO";
    CCU2D add_143_13 (.A0(cnt_delay[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt_delay[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n20502), .COUT(n20503), .S0(n2559[11]), 
          .S1(n2559[12]));   // g:/fpga/mxo2/system/project/oled12832.v(172[29:45])
    defparam add_143_13.INIT0 = 16'h5aaa;
    defparam add_143_13.INIT1 = 16'h5aaa;
    defparam add_143_13.INJECT1_0 = "NO";
    defparam add_143_13.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_127 (.A(cnt_init[0]), .B(n9817), .C(state_back[2]), 
         .D(n25755), .Z(n16_adj_5074)) /* synthesis lut_function=(!(A+!(B+(C (D))))) */ ;
    defparam i1_4_lut_adj_127.init = 16'h5444;
    LUT4 equal_1328_i11_2_lut_rep_357_3_lut_4_lut (.A(state[3]), .B(n25760), 
         .C(n25761), .D(state[0]), .Z(n25639)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(77[5:9])
    defparam equal_1328_i11_2_lut_rep_357_3_lut_4_lut.init = 16'hffef;
    CCU2D sub_1361_add_2_11 (.A0(cnt_delay[9]), .B0(num1_delay[9]), .C0(GND_net), 
          .D0(GND_net), .A1(cnt_delay[10]), .B1(num1_delay[10]), .C1(GND_net), 
          .D1(GND_net), .CIN(n20589), .COUT(n20590));
    defparam sub_1361_add_2_11.INIT0 = 16'h5999;
    defparam sub_1361_add_2_11.INIT1 = 16'h5999;
    defparam sub_1361_add_2_11.INJECT1_0 = "NO";
    defparam sub_1361_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_1361_add_2_9 (.A0(cnt_delay[7]), .B0(num1_delay[7]), .C0(GND_net), 
          .D0(GND_net), .A1(cnt_delay[8]), .B1(num1_delay[8]), .C1(GND_net), 
          .D1(GND_net), .CIN(n20588), .COUT(n20589));
    defparam sub_1361_add_2_9.INIT0 = 16'h5999;
    defparam sub_1361_add_2_9.INIT1 = 16'h5999;
    defparam sub_1361_add_2_9.INJECT1_0 = "NO";
    defparam sub_1361_add_2_9.INJECT1_1 = "NO";
    LUT4 cnt_scan_1__bdd_4_lut_22580 (.A(n25635), .B(num2[0]), .C(n25753), 
         .D(n25676), .Z(n25031)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+(C+!(D)))) */ ;
    defparam cnt_scan_1__bdd_4_lut_22580.init = 16'h8108;
    CCU2D sub_1361_add_2_7 (.A0(cnt_delay[5]), .B0(num1_delay[5]), .C0(GND_net), 
          .D0(GND_net), .A1(cnt_delay[6]), .B1(num1_delay[6]), .C1(GND_net), 
          .D1(GND_net), .CIN(n20587), .COUT(n20588));
    defparam sub_1361_add_2_7.INIT0 = 16'h5999;
    defparam sub_1361_add_2_7.INIT1 = 16'h5999;
    defparam sub_1361_add_2_7.INJECT1_0 = "NO";
    defparam sub_1361_add_2_7.INJECT1_1 = "NO";
    LUT4 n2421_bdd_4_lut_21993 (.A(cnt_scan[1]), .B(n25594), .C(num2[0]), 
         .D(n25753), .Z(n25030)) /* synthesis lut_function=(A (B (D))+!A !((C+!(D))+!B)) */ ;
    defparam n2421_bdd_4_lut_21993.init = 16'h8c00;
    LUT4 i1_3_lut_4_lut_adj_128 (.A(cnt_init[0]), .B(n25677), .C(n25650), 
         .D(num1_delay[3]), .Z(n4_adj_5104)) /* synthesis lut_function=(A ((C (D))+!B)+!A (C (D))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam i1_3_lut_4_lut_adj_128.init = 16'hf222;
    LUT4 i1_4_lut_adj_129 (.A(state[0]), .B(char[1]), .C(n16_adj_5105), 
         .D(n19_adj_5092), .Z(char_7__N_553[1])) /* synthesis lut_function=(A (B (D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_129.init = 16'hdc50;
    LUT4 i2_3_lut_4_lut_adj_130 (.A(state[3]), .B(n25760), .C(n10049), 
         .D(state[2]), .Z(n19_adj_5092)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(77[5:9])
    defparam i2_3_lut_4_lut_adj_130.init = 16'hfffe;
    PFUMX i59 (.BLUT(n28), .ALUT(n31_adj_5106), .C0(cnt_main[3]), .Z(n39));
    LUT4 i33_4_lut_adj_131 (.A(char[1]), .B(char_7__N_756[1]), .C(state[1]), 
         .D(n25646), .Z(n16_adj_5105)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam i33_4_lut_adj_131.init = 16'h0aca;
    LUT4 i1_4_lut_adj_132 (.A(n16111), .B(char[1]), .C(n4_adj_5107), .D(n36), 
         .Z(char_7__N_756[1])) /* synthesis lut_function=((B (C+(D))+!B (C))+!A) */ ;
    defparam i1_4_lut_adj_132.init = 16'hfdf5;
    FD1P3IX cnt_init_i0_i2 (.D(n1[2]), .SP(clk_c_enable_1359), .CD(n12024), 
            .CK(clk_c), .Q(cnt_init[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam cnt_init_i0_i2.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_339 (.A(num1[0]), .B(n1359), .Z(n25621)) /* synthesis lut_function=(A (B)) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(111[7] 142[14])
    defparam i1_2_lut_rep_339.init = 16'h8888;
    LUT4 i5918_4_lut_4_lut (.A(n25601), .B(n23698), .C(n30), .D(num2[0]), 
         .Z(n8725)) /* synthesis lut_function=(A (B (D))+!A (C)) */ ;
    defparam i5918_4_lut_4_lut.init = 16'hd850;
    LUT4 cnt_main_1__bdd_4_lut_22235 (.A(cnt_main[1]), .B(cnt_main[3]), 
         .C(cnt_main[0]), .D(cnt_main[2]), .Z(n58)) /* synthesis lut_function=(!(A (B (C (D)))+!A !(B+(C+(D))))) */ ;
    defparam cnt_main_1__bdd_4_lut_22235.init = 16'h7ffe;
    CCU2D sub_1361_add_2_5 (.A0(cnt_delay[3]), .B0(num1_delay[3]), .C0(GND_net), 
          .D0(GND_net), .A1(cnt_delay[4]), .B1(num1_delay[4]), .C1(GND_net), 
          .D1(GND_net), .CIN(n20586), .COUT(n20587));
    defparam sub_1361_add_2_5.INIT0 = 16'h5999;
    defparam sub_1361_add_2_5.INIT1 = 16'h5999;
    defparam sub_1361_add_2_5.INJECT1_0 = "NO";
    defparam sub_1361_add_2_5.INJECT1_1 = "NO";
    LUT4 i21065_3_lut_4_lut_4_lut (.A(n25601), .B(n16722), .C(n25589), 
         .D(num2[0]), .Z(n23942)) /* synthesis lut_function=(!(A (B)+!A (C+(D)))) */ ;
    defparam i21065_3_lut_4_lut_4_lut.init = 16'h2227;
    LUT4 i1_2_lut_rep_330_3_lut_4_lut (.A(state[3]), .B(n25760), .C(n25761), 
         .D(state[0]), .Z(n25612)) /* synthesis lut_function=(!(A+(B+!((D)+!C)))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(77[5:9])
    defparam i1_2_lut_rep_330_3_lut_4_lut.init = 16'h1101;
    FD1P3IX cnt_init_i0_i3 (.D(n1[3]), .SP(clk_c_enable_1359), .CD(n12024), 
            .CK(clk_c), .Q(cnt_init[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam cnt_init_i0_i3.GSR = "ENABLED";
    PFUMX i21878 (.BLUT(n25123), .ALUT(n25122), .C0(cnt_main[0]), .Z(n25124));
    LUT4 i9202_2_lut_3_lut_4_lut (.A(state[3]), .B(n25760), .C(clk_c_enable_1401), 
         .D(n8), .Z(n12017)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(77[5:9])
    defparam i9202_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i1_4_lut_adj_133 (.A(state[0]), .B(char[2]), .C(n16_adj_5108), 
         .D(n19_adj_5092), .Z(char_7__N_553[2])) /* synthesis lut_function=(A (B (D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_133.init = 16'hdc50;
    LUT4 i21068_3_lut_4_lut_4_lut (.A(n25601), .B(n24961), .C(n25594), 
         .D(num2[0]), .Z(n23945)) /* synthesis lut_function=(A (B)+!A (C (D))) */ ;
    defparam i21068_3_lut_4_lut_4_lut.init = 16'hd888;
    LUT4 i33_4_lut_adj_134 (.A(char[2]), .B(char_7__N_756[2]), .C(state[1]), 
         .D(n25646), .Z(n16_adj_5108)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam i33_4_lut_adj_134.init = 16'h0aca;
    LUT4 i21069_3_lut_3_lut_4_lut_4_lut (.A(n25601), .B(n23761), .C(n25594), 
         .D(num2[0]), .Z(n23946)) /* synthesis lut_function=(!(A (B)+!A ((D)+!C))) */ ;
    defparam i21069_3_lut_3_lut_4_lut_4_lut.init = 16'h2272;
    FD1P3IX cnt_init_i0_i4 (.D(n1[4]), .SP(clk_c_enable_1359), .CD(n12024), 
            .CK(clk_c), .Q(cnt_init[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam cnt_init_i0_i4.GSR = "ENABLED";
    PFUMX i21875 (.BLUT(n25120), .ALUT(n25119), .C0(cnt_scan[0]), .Z(n25121));
    LUT4 mux_414_Mux_23_i15_4_lut (.A(n25590), .B(n25624), .C(n25635), 
         .D(n25753), .Z(n16722)) /* synthesis lut_function=(A (((D)+!C)+!B)+!A (B (C (D))+!B (C))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(139[72:96])
    defparam mux_414_Mux_23_i15_4_lut.init = 16'hfa3a;
    LUT4 i1_3_lut_adj_135 (.A(char[2]), .B(cnt_main[4]), .C(n65), .Z(n41_adj_5109)) /* synthesis lut_function=(A (B+(C))) */ ;
    defparam i1_3_lut_adj_135.init = 16'ha8a8;
    PFUMX i21645 (.BLUT(n24682), .ALUT(n24681), .C0(cnt_scan[2]), .Z(n24683));
    CCU2D sub_1361_add_2_3 (.A0(cnt_delay[1]), .B0(num1_delay[1]), .C0(GND_net), 
          .D0(GND_net), .A1(cnt_delay[2]), .B1(num1_delay[2]), .C1(GND_net), 
          .D1(GND_net), .CIN(n20585), .COUT(n20586));
    defparam sub_1361_add_2_3.INIT0 = 16'h5999;
    defparam sub_1361_add_2_3.INIT1 = 16'h5999;
    defparam sub_1361_add_2_3.INJECT1_0 = "NO";
    defparam sub_1361_add_2_3.INJECT1_1 = "NO";
    FD1P3IX state_i0_i5 (.D(n32_adj_5065), .SP(clk_c_enable_1374), .CD(n16664), 
            .CK(clk_c), .Q(state[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam state_i0_i5.GSR = "ENABLED";
    FD1P3IX cnt_write_i0_i1 (.D(n2535[1]), .SP(clk_c_enable_1436), .CD(n12019), 
            .CK(clk_c), .Q(cnt_write[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam cnt_write_i0_i1.GSR = "ENABLED";
    CCU2D sub_1361_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt_delay[0]), .B1(num1_delay[0]), .C1(GND_net), 
          .D1(GND_net), .COUT(n20585));
    defparam sub_1361_add_2_1.INIT0 = 16'h0000;
    defparam sub_1361_add_2_1.INIT1 = 16'h5999;
    defparam sub_1361_add_2_1.INJECT1_0 = "NO";
    defparam sub_1361_add_2_1.INJECT1_1 = "NO";
    FD1P3IX cnt_write_i0_i2 (.D(n2535[2]), .SP(clk_c_enable_1436), .CD(n12019), 
            .CK(clk_c), .Q(cnt_write[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam cnt_write_i0_i2.GSR = "ENABLED";
    FD1P3IX cnt_write_i0_i3 (.D(n2535[3]), .SP(clk_c_enable_1436), .CD(n12019), 
            .CK(clk_c), .Q(cnt_write[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam cnt_write_i0_i3.GSR = "ENABLED";
    CCU2D add_143_11 (.A0(cnt_delay[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt_delay[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n20501), .COUT(n20502), .S0(n2559[9]), .S1(n2559[10]));   // g:/fpga/mxo2/system/project/oled12832.v(172[29:45])
    defparam add_143_11.INIT0 = 16'h5aaa;
    defparam add_143_11.INIT1 = 16'h5aaa;
    defparam add_143_11.INJECT1_0 = "NO";
    defparam add_143_11.INJECT1_1 = "NO";
    LUT4 i13350_2_lut_3_lut_4_lut_4_lut (.A(n25761), .B(state[0]), .C(n25760), 
         .D(state[3]), .Z(n5817[0])) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i13350_2_lut_3_lut_4_lut_4_lut.init = 16'h0008;
    LUT4 n25034_bdd_3_lut (.A(n25034), .B(n25031), .C(cnt_scan[1]), .Z(n25035)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25034_bdd_3_lut.init = 16'hcaca;
    LUT4 i21594_2_lut_rep_286_3_lut_4_lut_4_lut_4_lut (.A(n25761), .B(n25683), 
         .C(n25605), .D(n25684), .Z(clk_c_enable_1452)) /* synthesis lut_function=(!(A (B (C (D))+!B (C+!(D)))+!A (B (C)+!B (C+!(D))))) */ ;
    defparam i21594_2_lut_rep_286_3_lut_4_lut_4_lut_4_lut.init = 16'h0f8c;
    FD1P3IX state_i0_i4 (.D(n32_adj_5069), .SP(clk_c_enable_1374), .CD(n16664), 
            .CK(clk_c), .Q(state[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam state_i0_i4.GSR = "ENABLED";
    LUT4 i3438_2_lut_rep_340 (.A(n1359), .B(n1358), .Z(n25622)) /* synthesis lut_function=(!((B)+!A)) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(129[51:75])
    defparam i3438_2_lut_rep_340.init = 16'h2222;
    LUT4 i87_4_lut (.A(n25651), .B(n25677), .C(cnt_init[0]), .D(oled_dcn_N_888), 
         .Z(n79)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B)) */ ;
    defparam i87_4_lut.init = 16'hc4cc;
    LUT4 i1_4_lut_adj_136 (.A(state[0]), .B(char[3]), .C(n16_adj_5110), 
         .D(n19_adj_5092), .Z(char_7__N_553[3])) /* synthesis lut_function=(A (B (D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_136.init = 16'hdc50;
    LUT4 i21423_2_lut_rep_285_3_lut_4_lut_4_lut_4_lut (.A(n25761), .B(n25683), 
         .C(n25604), .D(n25684), .Z(clk_c_enable_1436)) /* synthesis lut_function=(!(A (B (C (D))+!B (C+!(D)))+!A (B (C)+!B (C+!(D))))) */ ;
    defparam i21423_2_lut_rep_285_3_lut_4_lut_4_lut_4_lut.init = 16'h0f8c;
    LUT4 n93_bdd_3_lut_22079_4_lut (.A(n1359), .B(n1358), .C(num1[0]), 
         .D(n1357), .Z(n25062)) /* synthesis lut_function=(!((B+!(C (D)+!C !(D)))+!A)) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(129[51:75])
    defparam n93_bdd_3_lut_22079_4_lut.init = 16'h2002;
    LUT4 mux_414_Mux_15_i15_4_lut_4_lut_4_lut (.A(n25667), .B(n25561), .C(n25676), 
         .D(n25601), .Z(n15_adj_5111)) /* synthesis lut_function=(!(A ((D)+!B)+!A !(B (C+!(D))+!B (C (D))))) */ ;
    defparam mux_414_Mux_15_i15_4_lut_4_lut_4_lut.init = 16'h50cc;
    LUT4 i33_4_lut_adj_137 (.A(char[3]), .B(char_7__N_756[3]), .C(state[1]), 
         .D(n25646), .Z(n16_adj_5110)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam i33_4_lut_adj_137.init = 16'h0aca;
    LUT4 i21081_3_lut_3_lut_4_lut_4_lut (.A(n25601), .B(n15_adj_5112), .C(n25594), 
         .D(num2[0]), .Z(n23958)) /* synthesis lut_function=(A (B)+!A !((D)+!C)) */ ;
    defparam i21081_3_lut_3_lut_4_lut_4_lut.init = 16'h88d8;
    LUT4 i2_3_lut_adj_138 (.A(cnt_main[0]), .B(n4_adj_5113), .C(n59), 
         .Z(char_7__N_756[3])) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;
    defparam i2_3_lut_adj_138.init = 16'hdcdc;
    LUT4 i21333_2_lut (.A(n3264), .B(n24047), .Z(clk_c_enable_1429)) /* synthesis lut_function=(A (B)) */ ;
    defparam i21333_2_lut.init = 16'h8888;
    CCU2D add_143_9 (.A0(cnt_delay[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt_delay[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n20500), .COUT(n20501), .S0(n2559[7]), .S1(n2559[8]));   // g:/fpga/mxo2/system/project/oled12832.v(172[29:45])
    defparam add_143_9.INIT0 = 16'h5aaa;
    defparam add_143_9.INIT1 = 16'h5aaa;
    defparam add_143_9.INJECT1_0 = "NO";
    defparam add_143_9.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_139 (.A(cnt_main[0]), .B(cnt_main[3]), .C(n24715), 
         .D(n24697), .Z(n68_adj_5114)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A !(B+!(D))) */ ;
    defparam i1_4_lut_adj_139.init = 16'hb3a0;
    LUT4 i1_2_lut_4_lut_adj_140 (.A(n25579), .B(n1355), .C(n1357), .D(n23306), 
         .Z(n23307)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(129[51:75])
    defparam i1_2_lut_4_lut_adj_140.init = 16'h2000;
    LUT4 i21332_4_lut (.A(n4432), .B(n4_adj_5115), .C(n25609), .D(n4434), 
         .Z(n24047)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B+!(C (D))))) */ ;
    defparam i21332_4_lut.init = 16'h3a0a;
    LUT4 mux_1117_i1_4_lut (.A(n4432), .B(n4434), .C(n25609), .D(n4_adj_5116), 
         .Z(n3189[0])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(41[4] 175[11])
    defparam mux_1117_i1_4_lut.init = 16'hca0a;
    LUT4 i1_4_lut_adj_141 (.A(state[0]), .B(char[4]), .C(n16_adj_5117), 
         .D(n19_adj_5092), .Z(char_7__N_553[4])) /* synthesis lut_function=(A (B (D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_141.init = 16'hdc50;
    LUT4 i33_4_lut_adj_142 (.A(char[4]), .B(n74), .C(state[1]), .D(n25646), 
         .Z(n16_adj_5117)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (B+((D)+!C)))) */ ;
    defparam i33_4_lut_adj_142.init = 16'h0a3a;
    LUT4 i1_4_lut_adj_143 (.A(n16111), .B(n89_adj_5118), .C(char[4]), 
         .D(n24915), .Z(n74)) /* synthesis lut_function=(A (B+!(C+!(D)))) */ ;
    defparam i1_4_lut_adj_143.init = 16'h8a88;
    CCU2D add_143_7 (.A0(cnt_delay[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt_delay[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n20499), .COUT(n20500), .S0(n2559[5]), .S1(n2559[6]));   // g:/fpga/mxo2/system/project/oled12832.v(172[29:45])
    defparam add_143_7.INIT0 = 16'h5aaa;
    defparam add_143_7.INIT1 = 16'h5aaa;
    defparam add_143_7.INJECT1_0 = "NO";
    defparam add_143_7.INJECT1_1 = "NO";
    PFUMX i133 (.BLUT(n76), .ALUT(n86), .C0(cnt_main[3]), .Z(n136));
    CCU2D add_143_5 (.A0(cnt_delay[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt_delay[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n20498), .COUT(n20499), .S0(n2559[3]), .S1(n2559[4]));   // g:/fpga/mxo2/system/project/oled12832.v(172[29:45])
    defparam add_143_5.INIT0 = 16'h5aaa;
    defparam add_143_5.INIT1 = 16'h5aaa;
    defparam add_143_5.INJECT1_0 = "NO";
    defparam add_143_5.INJECT1_1 = "NO";
    LUT4 mux_414_Mux_24_i15_4_lut (.A(num2[0]), .B(n14_adj_5119), .C(n25635), 
         .D(n25632), .Z(n15_adj_5120)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(139[72:96])
    defparam mux_414_Mux_24_i15_4_lut.init = 16'hcac0;
    LUT4 i1_3_lut_adj_144 (.A(cnt_main[0]), .B(n136), .C(n96), .Z(n105)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i1_3_lut_adj_144.init = 16'hecec;
    LUT4 i1_4_lut_adj_145 (.A(cnt_main[3]), .B(cnt_main[2]), .C(\tamp_data[3] ), 
         .D(time_data[9]), .Z(n96)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A ((D)+!B))) */ ;
    defparam i1_4_lut_adj_145.init = 16'h0ace;
    LUT4 n25047_bdd_3_lut_3_lut (.A(n25601), .B(n25044), .C(n25047), .Z(n25048)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam n25047_bdd_3_lut_3_lut.init = 16'he4e4;
    LUT4 i21077_3_lut_4_lut_4_lut (.A(n25601), .B(n23507), .C(n25589), 
         .D(num2[0]), .Z(n23954)) /* synthesis lut_function=(!(A (B)+!A (C+(D)))) */ ;
    defparam i21077_3_lut_4_lut_4_lut.init = 16'h2227;
    LUT4 i1_4_lut_adj_146 (.A(state[0]), .B(char[5]), .C(n16_adj_5121), 
         .D(n19_adj_5092), .Z(char_7__N_553[5])) /* synthesis lut_function=(A (B (D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_146.init = 16'hdc50;
    FD1P3IX cnt_write_i0_i4 (.D(n2535[4]), .SP(clk_c_enable_1436), .CD(n12019), 
            .CK(clk_c), .Q(cnt_write[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam cnt_write_i0_i4.GSR = "ENABLED";
    LUT4 i33_4_lut_adj_147 (.A(char[5]), .B(char_7__N_756[5]), .C(state[1]), 
         .D(n25646), .Z(n16_adj_5121)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam i33_4_lut_adj_147.init = 16'h0aca;
    FD1P3IX state_i0_i3 (.D(n21577), .SP(clk_c_enable_1374), .CD(n12116), 
            .CK(clk_c), .Q(state[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam state_i0_i3.GSR = "ENABLED";
    FD1P3IX state_i0_i2 (.D(n21575), .SP(clk_c_enable_1374), .CD(n12116), 
            .CK(clk_c), .Q(state[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam state_i0_i2.GSR = "ENABLED";
    FD1P3IX cnt_i0_i15 (.D(n167[15]), .SP(clk_c_enable_1401), .CD(n12017), 
            .CK(clk_c), .Q(cnt_c[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam cnt_i0_i15.GSR = "ENABLED";
    FD1P3AX state_i0_i1 (.D(n26497), .SP(clk_c_enable_1374), .CK(clk_c), 
            .Q(state[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam state_i0_i1.GSR = "ENABLED";
    FD1P3IX cnt_i0_i14 (.D(n167[14]), .SP(clk_c_enable_1401), .CD(n12017), 
            .CK(clk_c), .Q(cnt_c[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam cnt_i0_i14.GSR = "ENABLED";
    FD1P3IX cnt_i0_i13 (.D(n167[13]), .SP(clk_c_enable_1401), .CD(n12017), 
            .CK(clk_c), .Q(cnt_c[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam cnt_i0_i13.GSR = "ENABLED";
    FD1P3IX cnt_i0_i12 (.D(n167[12]), .SP(clk_c_enable_1401), .CD(n12017), 
            .CK(clk_c), .Q(cnt_c[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam cnt_i0_i12.GSR = "ENABLED";
    FD1P3IX cnt_i0_i0 (.D(n167[0]), .SP(clk_c_enable_1401), .CD(n12017), 
            .CK(clk_c), .Q(cnt[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam cnt_i0_i0.GSR = "ENABLED";
    LUT4 i1_3_lut_4_lut_adj_148 (.A(n25570), .B(n25755), .C(num1_delay[5]), 
         .D(cnt_init[0]), .Z(n16_adj_5122)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;
    defparam i1_3_lut_4_lut_adj_148.init = 16'h00e0;
    FD1P3IX cnt_i0_i11 (.D(n167[11]), .SP(clk_c_enable_1401), .CD(n12017), 
            .CK(clk_c), .Q(cnt_c[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam cnt_i0_i11.GSR = "ENABLED";
    FD1P3IX cnt_i0_i10 (.D(n167[10]), .SP(clk_c_enable_1401), .CD(n12017), 
            .CK(clk_c), .Q(cnt_c[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam cnt_i0_i10.GSR = "ENABLED";
    FD1P3IX cnt_i0_i9 (.D(n167[9]), .SP(clk_c_enable_1401), .CD(n12017), 
            .CK(clk_c), .Q(cnt_c[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam cnt_i0_i9.GSR = "ENABLED";
    FD1P3IX cnt_i0_i8 (.D(n167[8]), .SP(clk_c_enable_1401), .CD(n12017), 
            .CK(clk_c), .Q(cnt_c[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam cnt_i0_i8.GSR = "ENABLED";
    FD1P3IX cnt_i0_i7 (.D(n167[7]), .SP(clk_c_enable_1401), .CD(n12017), 
            .CK(clk_c), .Q(cnt_c[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam cnt_i0_i7.GSR = "ENABLED";
    FD1P3IX cnt_i0_i6 (.D(n167[6]), .SP(clk_c_enable_1401), .CD(n12017), 
            .CK(clk_c), .Q(cnt_c[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam cnt_i0_i6.GSR = "ENABLED";
    FD1P3IX cnt_i0_i5 (.D(n167[5]), .SP(clk_c_enable_1401), .CD(n12017), 
            .CK(clk_c), .Q(cnt_c[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam cnt_i0_i5.GSR = "ENABLED";
    FD1P3IX cnt_i0_i4 (.D(n167[4]), .SP(clk_c_enable_1401), .CD(n12017), 
            .CK(clk_c), .Q(cnt[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam cnt_i0_i4.GSR = "ENABLED";
    FD1P3IX cnt_i0_i3 (.D(n167[3]), .SP(clk_c_enable_1401), .CD(n12017), 
            .CK(clk_c), .Q(cnt[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam cnt_i0_i3.GSR = "ENABLED";
    PFUMX i21848 (.BLUT(n25062), .ALUT(n93), .C0(n1356), .Z(n25063));
    LUT4 i1_4_lut_adj_149 (.A(char[5]), .B(n25124), .C(n9), .D(n15942), 
         .Z(char_7__N_756[5])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((D)+!B)) */ ;
    defparam i1_4_lut_adj_149.init = 16'ha0ec;
    FD1P3IX cnt_i0_i2 (.D(n167[2]), .SP(clk_c_enable_1401), .CD(n12017), 
            .CK(clk_c), .Q(cnt[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam cnt_i0_i2.GSR = "ENABLED";
    LUT4 unary_minus_2211_inv_0_i1_1_lut_rep_403 (.A(num1[0]), .Z(n25685)) /* synthesis lut_function=(!(A)) */ ;
    defparam unary_minus_2211_inv_0_i1_1_lut_rep_403.init = 16'h5555;
    LUT4 i1_4_lut_adj_150 (.A(state[0]), .B(char[6]), .C(n16_adj_5123), 
         .D(n19_adj_5092), .Z(char_7__N_553[6])) /* synthesis lut_function=(A (B (D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_150.init = 16'hdc50;
    LUT4 i18413_1_lut (.A(n3599), .Z(n21240)) /* synthesis lut_function=(!(A)) */ ;
    defparam i18413_1_lut.init = 16'h5555;
    LUT4 i1_3_lut_4_lut_adj_151 (.A(n25570), .B(n25755), .C(num1_delay[8]), 
         .D(cnt_init[0]), .Z(n16_adj_5124)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;
    defparam i1_3_lut_4_lut_adj_151.init = 16'h00e0;
    LUT4 i33_4_lut_adj_152 (.A(char[6]), .B(char_7__N_756[6]), .C(state[1]), 
         .D(n25646), .Z(n16_adj_5123)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam i33_4_lut_adj_152.init = 16'h0aca;
    LUT4 mux_415_Mux_22_i92_3_lut_4_lut_3_lut (.A(num1[0]), .B(n1358), .C(n1359), 
         .Z(n92)) /* synthesis lut_function=(A (B (C))+!A !(B)) */ ;
    defparam mux_415_Mux_22_i92_3_lut_4_lut_3_lut.init = 16'h9191;
    LUT4 i2_4_lut_adj_153 (.A(n37_adj_5125), .B(cnt_main[0]), .C(n43_adj_5076), 
         .D(n25805), .Z(char_7__N_756[6])) /* synthesis lut_function=(A+(B (C)+!B (C+(D)))) */ ;
    defparam i2_4_lut_adj_153.init = 16'hfbfa;
    LUT4 i2_4_lut_adj_154 (.A(cnt_main[0]), .B(n15942), .C(n61), .D(n45), 
         .Z(n37_adj_5125)) /* synthesis lut_function=(!(A (B+!(C+(D)))+!A (B+!(C)))) */ ;
    defparam i2_4_lut_adj_154.init = 16'h3230;
    LUT4 i3042_1_lut (.A(cnt_write[0]), .Z(n4_adj_5126)) /* synthesis lut_function=(!(A)) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(147[7] 167[14])
    defparam i3042_1_lut.init = 16'h5555;
    PFUMX i21840 (.BLUT(n25046), .ALUT(n25045), .C0(cnt_scan[1]), .Z(n25047));
    LUT4 i1_3_lut_4_lut_adj_155 (.A(n25570), .B(n25755), .C(num1_delay[13]), 
         .D(cnt_init[0]), .Z(n16_adj_5127)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;
    defparam i1_3_lut_4_lut_adj_155.init = 16'h00e0;
    LUT4 i1_3_lut_4_lut_adj_156 (.A(n25570), .B(n25755), .C(num1_delay[14]), 
         .D(cnt_init[0]), .Z(n16_adj_5128)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;
    defparam i1_3_lut_4_lut_adj_156.init = 16'h00e0;
    LUT4 n93_bdd_4_lut_4_lut (.A(num1[0]), .B(n25622), .C(n1356), .D(n1357), 
         .Z(n25064)) /* synthesis lut_function=(!(A+!(B (C (D)+!C !(D))))) */ ;
    defparam n93_bdd_4_lut_4_lut.init = 16'h4004;
    CCU2D add_143_3 (.A0(cnt_delay[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt_delay[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n20497), .COUT(n20498), .S0(n2559[1]), .S1(n2559[2]));   // g:/fpga/mxo2/system/project/oled12832.v(172[29:45])
    defparam add_143_3.INIT0 = 16'h5aaa;
    defparam add_143_3.INIT1 = 16'h5aaa;
    defparam add_143_3.INJECT1_0 = "NO";
    defparam add_143_3.INJECT1_1 = "NO";
    LUT4 mux_415_Mux_30_i92_3_lut_rep_317_4_lut_4_lut_3_lut (.A(num1[0]), 
         .B(n1358), .C(n1359), .Z(n25599)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B+!(C)))) */ ;
    defparam mux_415_Mux_30_i92_3_lut_rep_317_4_lut_4_lut_3_lut.init = 16'h1818;
    LUT4 n20924_bdd_4_lut_21839 (.A(n25753), .B(cnt_scan[1]), .C(num2[0]), 
         .D(n25594), .Z(n25044)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C (D)))+!A !(B (C (D))+!B !(C+!(D))))) */ ;
    defparam n20924_bdd_4_lut_21839.init = 16'h6900;
    LUT4 i1_2_lut_4_lut_4_lut (.A(num1[0]), .B(n25566), .C(n25622), .D(cnt_scan[0]), 
         .Z(n23360)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_2_lut_4_lut_4_lut.init = 16'h4000;
    LUT4 i1_2_lut_3_lut_3_lut (.A(num1[0]), .B(n1358), .C(n1359), .Z(n23306)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_3_lut.init = 16'h1010;
    LUT4 n26417_bdd_4_lut (.A(n26417), .B(n26416), .C(n25601), .D(num2[0]), 
         .Z(n26778)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam n26417_bdd_4_lut.init = 16'hca00;
    LUT4 n92_bdd_4_lut_4_lut (.A(num1[0]), .B(n1358), .C(n1356), .D(n1359), 
         .Z(n24905)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C+!(D)))+!A (B ((D)+!C)+!B !(D)))) */ ;
    defparam n92_bdd_4_lut_4_lut.init = 16'h13c0;
    LUT4 mux_131_Mux_2_i11_4_lut_4_lut (.A(num1[0]), .B(n25557), .C(cnt_scan[0]), 
         .D(n863), .Z(n11_adj_5129)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (C+!(D)))) */ ;
    defparam mux_131_Mux_2_i11_4_lut_4_lut.init = 16'h2f20;
    LUT4 i2_4_lut_adj_157 (.A(n11_adj_5073), .B(n25719), .C(n21240), .D(cnt_scan[2]), 
         .Z(n21243)) /* synthesis lut_function=(!(A+(B ((D)+!C)+!B !(C (D))))) */ ;
    defparam i2_4_lut_adj_157.init = 16'h1040;
    LUT4 i1_3_lut_3_lut (.A(num1[0]), .B(n1358), .C(n1359), .Z(n23415)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i1_3_lut_3_lut.init = 16'hf7f7;
    LUT4 n23900_bdd_4_lut_4_lut (.A(cnt_scan[0]), .B(cnt_scan[3]), .C(n29_adj_5066), 
         .D(n16_adj_5130), .Z(n25037)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;
    defparam n23900_bdd_4_lut_4_lut.init = 16'hd1c0;
    LUT4 i21236_4_lut_4_lut (.A(cnt_scan[0]), .B(n23869), .C(n25412), 
         .D(n62), .Z(n11_adj_5131)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;
    defparam i21236_4_lut_4_lut.init = 16'hf4b0;
    LUT4 i1_4_lut_adj_158 (.A(state[0]), .B(num1_delay[1]), .C(n16_adj_5132), 
         .D(n27_adj_5133), .Z(num1_delay_15__N_605[1])) /* synthesis lut_function=(A (B (D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_158.init = 16'hdc50;
    LUT4 i33_4_lut_adj_159 (.A(num1_delay[1]), .B(num1_delay_15__N_780[1]), 
         .C(state[2]), .D(n16443), .Z(n16_adj_5132)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam i33_4_lut_adj_159.init = 16'h0aca;
    LUT4 i1_4_lut_adj_160 (.A(cnt_init[0]), .B(num1_delay[1]), .C(n25559), 
         .D(n25650), .Z(num1_delay_15__N_780[1])) /* synthesis lut_function=(A (B (D))+!A (B (C+(D)))) */ ;
    defparam i1_4_lut_adj_160.init = 16'hcc40;
    LUT4 mux_1283_i1_4_lut_3_lut (.A(cnt_scan[0]), .B(n3599), .C(n322), 
         .Z(cnt_scan_4__N_682[0])) /* synthesis lut_function=(A (B (C))+!A !(B)) */ ;
    defparam mux_1283_i1_4_lut_3_lut.init = 16'h9191;
    LUT4 cnt_scan_2__bdd_3_lut_21644 (.A(x_ph[3]), .B(cnt_scan[0]), .C(cnt_scan[1]), 
         .Z(n24681)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;
    defparam cnt_scan_2__bdd_3_lut_21644.init = 16'h0202;
    LUT4 i21462_4_lut (.A(state[0]), .B(num1_delay[2]), .C(n16726), .D(n27_adj_5133), 
         .Z(num1_delay_15__N_605[2])) /* synthesis lut_function=(A (B+!(D))+!A (B (C)+!B !((D)+!C))) */ ;
    defparam i21462_4_lut.init = 16'hc8fa;
    LUT4 i41_4_lut (.A(num1_delay[2]), .B(n16443), .C(state[2]), .D(n23209), 
         .Z(n16726)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;
    defparam i41_4_lut.init = 16'hfaca;
    LUT4 i1_4_lut_adj_161 (.A(cnt_init[0]), .B(num1_delay[2]), .C(n15_adj_5134), 
         .D(n25650), .Z(n23209)) /* synthesis lut_function=(A (B (D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_161.init = 16'hdc50;
    LUT4 i1_4_lut_adj_162 (.A(num1_delay[2]), .B(n25755), .C(n25651), 
         .D(oled_dcn_N_888), .Z(n15_adj_5134)) /* synthesis lut_function=(A (B+(C))+!A !((D)+!C)) */ ;
    defparam i1_4_lut_adj_162.init = 16'ha8f8;
    LUT4 i2_3_lut_3_lut (.A(cnt_scan[0]), .B(n25566), .C(n25599), .Z(n16_adj_5085)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i2_3_lut_3_lut.init = 16'h4040;
    LUT4 i1_4_lut_adj_163 (.A(state[0]), .B(num1_delay[3]), .C(n16_adj_5135), 
         .D(n27_adj_5133), .Z(num1_delay_15__N_605[3])) /* synthesis lut_function=(A (B (D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_163.init = 16'hdc50;
    LUT4 i33_4_lut_adj_164 (.A(num1_delay[3]), .B(num1_delay_15__N_780[3]), 
         .C(state[2]), .D(n16443), .Z(n16_adj_5135)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam i33_4_lut_adj_164.init = 16'h0aca;
    LUT4 i2_4_lut_adj_165 (.A(cnt_init[0]), .B(n4_adj_5104), .C(num1_delay[3]), 
         .D(n25559), .Z(num1_delay_15__N_780[3])) /* synthesis lut_function=(A (B)+!A (B+(C (D)))) */ ;
    defparam i2_4_lut_adj_165.init = 16'hdccc;
    LUT4 i1_3_lut_3_lut_adj_166 (.A(cnt_scan[0]), .B(x_pl[5]), .C(cnt_scan[1]), 
         .Z(n23099)) /* synthesis lut_function=((B (C))+!A) */ ;
    defparam i1_3_lut_3_lut_adj_166.init = 16'hd5d5;
    LUT4 i1_2_lut_2_lut (.A(cnt_scan[0]), .B(num2[0]), .Z(n23422)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i1_2_lut_2_lut.init = 16'hdddd;
    LUT4 i13537_2_lut_2_lut (.A(cnt_scan[0]), .B(n1423), .Z(n16_adj_5136)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i13537_2_lut_2_lut.init = 16'h4444;
    LUT4 n1354_bdd_4_lut_22276 (.A(n25599), .B(n1357), .C(n1356), .D(n25622), 
         .Z(n25060)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A ((C+!(D))+!B))) */ ;
    defparam n1354_bdd_4_lut_22276.init = 16'h2c20;
    LUT4 i9301_2_lut_3_lut (.A(n25605), .B(n2557), .C(state[0]), .Z(n12116)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i9301_2_lut_3_lut.init = 16'he0e0;
    PFUMX i21835 (.BLUT(n23900), .ALUT(n25037), .C0(cnt_scan[4]), .Z(n25038));
    LUT4 i1_4_lut_adj_167 (.A(state[0]), .B(num1_delay[4]), .C(n16_adj_5137), 
         .D(n27_adj_5133), .Z(num1_delay_15__N_605[4])) /* synthesis lut_function=(A (B (D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_167.init = 16'hdc50;
    LUT4 i33_4_lut_adj_168 (.A(num1_delay[4]), .B(num1_delay_15__N_780[4]), 
         .C(state[2]), .D(n16443), .Z(n16_adj_5137)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam i33_4_lut_adj_168.init = 16'h0aca;
    LUT4 i1_4_lut_adj_169 (.A(cnt_init[0]), .B(num1_delay[4]), .C(n25559), 
         .D(n25650), .Z(num1_delay_15__N_780[4])) /* synthesis lut_function=(A (B (D))+!A (B (C+(D)))) */ ;
    defparam i1_4_lut_adj_169.init = 16'hcc40;
    LUT4 i13351_2_lut_2_lut (.A(cnt_scan[0]), .B(n1425), .Z(n16_adj_5138)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i13351_2_lut_2_lut.init = 16'h4444;
    LUT4 i17787_2_lut_3_lut_3_lut (.A(cnt_scan[0]), .B(n25557), .C(num1[0]), 
         .Z(n8_adj_5139)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;
    defparam i17787_2_lut_3_lut_3_lut.init = 16'h0202;
    LUT4 n1058_bdd_2_lut_21953_2_lut (.A(cnt_scan[0]), .B(n25214), .Z(n25215)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam n1058_bdd_2_lut_21953_2_lut.init = 16'h4444;
    LUT4 i1_4_lut_adj_170 (.A(state[0]), .B(num1_delay[5]), .C(n16_adj_5140), 
         .D(n27_adj_5133), .Z(num1_delay_15__N_605[5])) /* synthesis lut_function=(A (B (D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_170.init = 16'hdc50;
    LUT4 i33_4_lut_adj_171 (.A(num1_delay[5]), .B(num1_delay_15__N_780[5]), 
         .C(state[2]), .D(n16443), .Z(n16_adj_5140)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam i33_4_lut_adj_171.init = 16'h0aca;
    LUT4 i1_4_lut_adj_172 (.A(n25620), .B(num1_delay[5]), .C(n16_adj_5122), 
         .D(n25650), .Z(num1_delay_15__N_780[5])) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_172.init = 16'hfefa;
    LUT4 i21273_3_lut_3_lut (.A(cnt_scan[0]), .B(n2030[29]), .C(n15_adj_5111), 
         .Z(n2162[21])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i21273_3_lut_3_lut.init = 16'he4e4;
    LUT4 i138_4_lut (.A(cnt_main[0]), .B(time_data[13]), .C(cnt_main[2]), 
         .D(time_data[21]), .Z(n76)) /* synthesis lut_function=(!(A (C+(D))+!A (B+!(C)))) */ ;
    defparam i138_4_lut.init = 16'h101a;
    LUT4 cnt_main_3__bdd_4_lut_22173 (.A(cnt_main[3]), .B(cnt_main[0]), 
         .C(cnt_main[1]), .D(cnt_main[2]), .Z(n25068)) /* synthesis lut_function=(!(A (C (D))+!A !(B (C)+!B (C+(D))))) */ ;
    defparam cnt_main_3__bdd_4_lut_22173.init = 16'h5bfa;
    LUT4 n20748_bdd_4_lut_4_lut (.A(cnt_scan[0]), .B(cnt_scan[2]), .C(n25048), 
         .D(n20748), .Z(n25186)) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)+!B (D)))) */ ;
    defparam n20748_bdd_4_lut_4_lut.init = 16'h7340;
    LUT4 n23282_bdd_4_lut (.A(n25645), .B(cnt_main[3]), .C(x_pl[5]), .D(cnt_main[1]), 
         .Z(n25073)) /* synthesis lut_function=(A (B (D)+!B !((D)+!C))+!A !(B+((D)+!C))) */ ;
    defparam n23282_bdd_4_lut.init = 16'h8830;
    LUT4 mux_3021_i1_4_lut (.A(n9), .B(n5817[0]), .C(n25587), .D(n16666), 
         .Z(n5820[0])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B+!(C))) */ ;
    defparam mux_3021_i1_4_lut.init = 16'hc5cf;
    LUT4 i21561_3_lut_3_lut_3_lut (.A(cnt_scan[0]), .B(n25601), .C(n25676), 
         .Z(n23861)) /* synthesis lut_function=(A+((C)+!B)) */ ;
    defparam i21561_3_lut_3_lut_3_lut.init = 16'hfbfb;
    LUT4 i1_4_lut_adj_173 (.A(state[0]), .B(num1_delay[6]), .C(n16_adj_5141), 
         .D(n27_adj_5133), .Z(num1_delay_15__N_605[6])) /* synthesis lut_function=(A (B (D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_173.init = 16'hdc50;
    LUT4 i1_2_lut_rep_404 (.A(cnt_scan[2]), .B(cnt_scan[1]), .Z(n25686)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_404.init = 16'heeee;
    LUT4 n20927_bdd_4_lut_21927 (.A(n25676), .B(n25601), .C(n25635), .D(n25753), 
         .Z(n25074)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A !(B (C (D))+!B !(C+(D))))) */ ;
    defparam n20927_bdd_4_lut_21927.init = 16'h4801;
    LUT4 i33_4_lut_adj_174 (.A(num1_delay[6]), .B(num1_delay_15__N_780[6]), 
         .C(state[2]), .D(n16443), .Z(n16_adj_5141)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam i33_4_lut_adj_174.init = 16'h0aca;
    LUT4 i1_4_lut_adj_175 (.A(cnt_init[0]), .B(num1_delay[6]), .C(n25559), 
         .D(n25650), .Z(num1_delay_15__N_780[6])) /* synthesis lut_function=(A (B (D))+!A (B (C+(D)))) */ ;
    defparam i1_4_lut_adj_175.init = 16'hcc40;
    LUT4 i1_2_lut_rep_332_3_lut_4_lut (.A(cnt_scan[2]), .B(cnt_scan[1]), 
         .C(cnt_scan[3]), .D(cnt_scan[0]), .Z(n25614)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;
    defparam i1_2_lut_rep_332_3_lut_4_lut.init = 16'hffef;
    LUT4 i1_2_lut_rep_378_3_lut (.A(cnt_scan[2]), .B(cnt_scan[1]), .C(cnt_scan[0]), 
         .Z(n25660)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_378_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_334_3_lut_4_lut (.A(cnt_scan[2]), .B(cnt_scan[1]), 
         .C(cnt_scan[3]), .D(cnt_scan[0]), .Z(n25616)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_2_lut_rep_334_3_lut_4_lut.init = 16'h0100;
    LUT4 i1_4_lut_adj_176 (.A(state[0]), .B(num1_delay[7]), .C(n16_adj_5142), 
         .D(n27_adj_5133), .Z(num1_delay_15__N_605[7])) /* synthesis lut_function=(A (B (D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_176.init = 16'hdc50;
    LUT4 cnt_scan_2__bdd_3_lut_21663 (.A(x_pl[3]), .B(cnt_scan[0]), .C(cnt_scan[1]), 
         .Z(n24682)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam cnt_scan_2__bdd_3_lut_21663.init = 16'h8080;
    LUT4 i4269_3_lut_3_lut_4_lut (.A(cnt_scan[2]), .B(cnt_scan[1]), .C(cnt_scan[3]), 
         .D(cnt_scan[0]), .Z(n8418)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !(C+!(D)))) */ ;
    defparam i4269_3_lut_3_lut_4_lut.init = 16'he1e0;
    LUT4 i2_4_lut_adj_177 (.A(\tamp_data[0] ), .B(n25672), .C(time_data[4]), 
         .D(cnt_main[1]), .Z(n31_adj_5106)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i2_4_lut_adj_177.init = 16'hc088;
    LUT4 i33_4_lut_adj_178 (.A(num1_delay[7]), .B(num1_delay_15__N_780[7]), 
         .C(state[2]), .D(n16443), .Z(n16_adj_5142)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam i33_4_lut_adj_178.init = 16'h0aca;
    LUT4 i2_4_lut_adj_179 (.A(cnt_init[0]), .B(n4_adj_5103), .C(num1_delay[7]), 
         .D(n25559), .Z(num1_delay_15__N_780[7])) /* synthesis lut_function=(A (B)+!A (B+(C (D)))) */ ;
    defparam i2_4_lut_adj_179.init = 16'hdccc;
    LUT4 mux_414_Mux_16_i15_4_lut_4_lut (.A(n25676), .B(n25635), .C(n25753), 
         .D(num2[0]), .Z(n15_adj_5143)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;
    defparam mux_414_Mux_16_i15_4_lut_4_lut.init = 16'hd1c0;
    LUT4 i1_4_lut_adj_180 (.A(state[0]), .B(num1_delay[8]), .C(n16_adj_5144), 
         .D(n27_adj_5133), .Z(num1_delay_15__N_605[8])) /* synthesis lut_function=(A (B (D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_180.init = 16'hdc50;
    PFUMX i21833 (.BLUT(n25035), .ALUT(n25030), .C0(n25574), .Z(n25036));
    LUT4 i33_4_lut_adj_181 (.A(num1_delay[8]), .B(num1_delay_15__N_780[8]), 
         .C(state[2]), .D(n16443), .Z(n16_adj_5144)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam i33_4_lut_adj_181.init = 16'h0aca;
    LUT4 i1_4_lut_adj_182 (.A(n25620), .B(num1_delay[8]), .C(n16_adj_5124), 
         .D(n25650), .Z(num1_delay_15__N_780[8])) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_182.init = 16'hfefa;
    LUT4 n20924_bdd_4_lut_4_lut (.A(n25676), .B(num2[0]), .C(n25635), 
         .D(n25753), .Z(n25046)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B (C+(D)))) */ ;
    defparam n20924_bdd_4_lut_4_lut.init = 16'h8069;
    LUT4 n2423_bdd_4_lut_4_lut (.A(n25676), .B(n25753), .C(num2[0]), .D(n25635), 
         .Z(n24961)) /* synthesis lut_function=(A (B (C (D))+!B !(C (D)+!C !(D)))+!A !(B (C+(D))+!B !(C))) */ ;
    defparam n2423_bdd_4_lut_4_lut.init = 16'h9234;
    FD1P3IX cnt_i0_i1 (.D(n167[1]), .SP(clk_c_enable_1401), .CD(n12017), 
            .CK(clk_c), .Q(cnt[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam cnt_i0_i1.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_183 (.A(state[0]), .B(num1_delay[9]), .C(n16_adj_5145), 
         .D(n27_adj_5133), .Z(num1_delay_15__N_605[9])) /* synthesis lut_function=(A (B (D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_183.init = 16'hdc50;
    LUT4 i33_4_lut_adj_184 (.A(num1_delay[9]), .B(num1_delay_15__N_780[9]), 
         .C(state[2]), .D(n16443), .Z(n16_adj_5145)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam i33_4_lut_adj_184.init = 16'h0aca;
    LUT4 i1_4_lut_adj_185 (.A(cnt_init[0]), .B(num1_delay[9]), .C(n25559), 
         .D(n25650), .Z(num1_delay_15__N_780[9])) /* synthesis lut_function=(A (B (D))+!A (B (C+(D)))) */ ;
    defparam i1_4_lut_adj_185.init = 16'hcc40;
    PFUMX i21831 (.BLUT(n25033), .ALUT(n25032), .C0(n25635), .Z(n25034));
    LUT4 i2_4_lut_adj_186 (.A(\tamp_data[8] ), .B(n25764), .C(\tamp_data[4] ), 
         .D(cnt_main[0]), .Z(n28)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i2_4_lut_adj_186.init = 16'hc088;
    LUT4 i1_4_lut_adj_187 (.A(state[0]), .B(num1_delay[10]), .C(n16_adj_5146), 
         .D(n27_adj_5133), .Z(num1_delay_15__N_605[10])) /* synthesis lut_function=(A (B (D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_187.init = 16'hdc50;
    LUT4 cnt_main_1__bdd_4_lut_22236 (.A(cnt_main[1]), .B(cnt_main[2]), 
         .C(cnt_main[3]), .D(cnt_main[4]), .Z(n16666)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B+((D)+!C))) */ ;
    defparam cnt_main_1__bdd_4_lut_22236.init = 16'hffe7;
    LUT4 i33_4_lut_adj_188 (.A(num1_delay[10]), .B(num1_delay_15__N_780[10]), 
         .C(state[2]), .D(n16443), .Z(n16_adj_5146)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam i33_4_lut_adj_188.init = 16'h0aca;
    LUT4 i1_4_lut_adj_189 (.A(cnt_init[0]), .B(num1_delay[10]), .C(n25559), 
         .D(n25650), .Z(num1_delay_15__N_780[10])) /* synthesis lut_function=(A (B (D))+!A (B (C+(D)))) */ ;
    defparam i1_4_lut_adj_189.init = 16'hcc40;
    LUT4 cnt_main_0__bdd_4_lut_21877 (.A(cnt_main[1]), .B(cnt_main[2]), 
         .C(time_data[22]), .D(time_data[10]), .Z(n25122)) /* synthesis lut_function=(!(A+!(B (D)+!B (C)))) */ ;
    defparam cnt_main_0__bdd_4_lut_21877.init = 16'h5410;
    LUT4 i1_4_lut_adj_190 (.A(state[0]), .B(num1_delay[11]), .C(n16_adj_5147), 
         .D(n27_adj_5133), .Z(num1_delay_15__N_605[11])) /* synthesis lut_function=(A (B (D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_190.init = 16'hdc50;
    LUT4 i33_4_lut_adj_191 (.A(num1_delay[11]), .B(num1_delay_15__N_780[11]), 
         .C(state[2]), .D(n16443), .Z(n16_adj_5147)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam i33_4_lut_adj_191.init = 16'h0aca;
    LUT4 cnt_main_0__bdd_4_lut_22353 (.A(cnt_main[1]), .B(cnt_main[2]), 
         .C(time_data[18]), .D(time_data[14]), .Z(n25123)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)))) */ ;
    defparam cnt_main_0__bdd_4_lut_22353.init = 16'h6420;
    LUT4 i1_4_lut_adj_192 (.A(cnt_init[0]), .B(num1_delay[11]), .C(n25559), 
         .D(n25650), .Z(num1_delay_15__N_780[11])) /* synthesis lut_function=(A (B (D))+!A (B (C+(D)))) */ ;
    defparam i1_4_lut_adj_192.init = 16'hcc40;
    LUT4 i17783_4_lut_4_lut_4_lut (.A(n25676), .B(n25753), .C(n4_adj_5148), 
         .D(n25601), .Z(n2030[29])) /* synthesis lut_function=(!(A (B (C+(D))+!B (C))+!A (C+!(D)))) */ ;
    defparam i17783_4_lut_4_lut_4_lut.init = 16'h070a;
    LUT4 i1_4_lut_adj_193 (.A(state[0]), .B(num1_delay[12]), .C(n16_adj_5149), 
         .D(n27_adj_5133), .Z(num1_delay_15__N_605[12])) /* synthesis lut_function=(A (B (D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_193.init = 16'hdc50;
    LUT4 i33_4_lut_adj_194 (.A(num1_delay[12]), .B(num1_delay_15__N_780[12]), 
         .C(state[2]), .D(n16443), .Z(n16_adj_5149)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam i33_4_lut_adj_194.init = 16'h0aca;
    LUT4 i1_4_lut_adj_195 (.A(cnt_init[0]), .B(num1_delay[12]), .C(n25559), 
         .D(n25650), .Z(num1_delay_15__N_780[12])) /* synthesis lut_function=(A (B (D))+!A (B (C+(D)))) */ ;
    defparam i1_4_lut_adj_195.init = 16'hcc40;
    LUT4 n20924_bdd_3_lut_4_lut (.A(n25676), .B(n25753), .C(num2[0]), 
         .D(n25635), .Z(n25045)) /* synthesis lut_function=(!((B+!(C (D)+!C !(D)))+!A)) */ ;
    defparam n20924_bdd_3_lut_4_lut.init = 16'h2002;
    LUT4 i17679_4_lut_4_lut_then_4_lut (.A(cnt_main[1]), .B(cnt_main[0]), 
         .C(cnt_main[4]), .D(cnt_main[2]), .Z(n25770)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(53[12:40])
    defparam i17679_4_lut_4_lut_then_4_lut.init = 16'h78f0;
    LUT4 i1_4_lut_adj_196 (.A(state[0]), .B(num1_delay[13]), .C(n16_adj_5150), 
         .D(n27_adj_5133), .Z(num1_delay_15__N_605[13])) /* synthesis lut_function=(A (B (D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_196.init = 16'hdc50;
    LUT4 i33_4_lut_adj_197 (.A(num1_delay[13]), .B(num1_delay_15__N_780[13]), 
         .C(state[2]), .D(n16443), .Z(n16_adj_5150)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam i33_4_lut_adj_197.init = 16'h0aca;
    LUT4 i1_4_lut_adj_198 (.A(n25620), .B(num1_delay[13]), .C(n16_adj_5127), 
         .D(n25650), .Z(num1_delay_15__N_780[13])) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_198.init = 16'hfefa;
    LUT4 cnt_scan_0__bdd_3_lut_4_lut (.A(n25676), .B(n25753), .C(num2[0]), 
         .D(n25635), .Z(n25369)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam cnt_scan_0__bdd_3_lut_4_lut.init = 16'h0002;
    LUT4 n26452_bdd_3_lut_4_lut (.A(n23942), .B(cnt_scan[2]), .C(cnt_scan[1]), 
         .D(n26451), .Z(n26453)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;
    defparam n26452_bdd_3_lut_4_lut.init = 16'hf808;
    LUT4 i1_4_lut_adj_199 (.A(state[0]), .B(num1_delay[14]), .C(n16_adj_5151), 
         .D(n27_adj_5133), .Z(num1_delay_15__N_605[14])) /* synthesis lut_function=(A (B (D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_199.init = 16'hdc50;
    LUT4 i33_4_lut_adj_200 (.A(num1_delay[14]), .B(num1_delay_15__N_780[14]), 
         .C(state[2]), .D(n16443), .Z(n16_adj_5151)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam i33_4_lut_adj_200.init = 16'h0aca;
    PFUMX i22167 (.BLUT(n25790), .ALUT(n25791), .C0(cnt_main[2]), .Z(num1_7__N_724[3]));
    LUT4 i1_4_lut_adj_201 (.A(n25620), .B(num1_delay[14]), .C(n16_adj_5128), 
         .D(n25650), .Z(num1_delay_15__N_780[14])) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_201.init = 16'hfefa;
    LUT4 i17679_4_lut_4_lut_else_4_lut (.A(cnt_main[4]), .Z(n25769)) /* synthesis lut_function=(A) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(53[12:40])
    defparam i17679_4_lut_4_lut_else_4_lut.init = 16'haaaa;
    LUT4 i1_4_lut_adj_202 (.A(state[0]), .B(num1_delay[15]), .C(n16_adj_5152), 
         .D(n27_adj_5133), .Z(num1_delay_15__N_605[15])) /* synthesis lut_function=(A (B (D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_202.init = 16'hdc50;
    LUT4 i33_4_lut_adj_203 (.A(num1_delay[15]), .B(num1_delay_15__N_780[15]), 
         .C(state[2]), .D(n16443), .Z(n16_adj_5152)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;
    defparam i33_4_lut_adj_203.init = 16'h0aca;
    LUT4 i1_4_lut_adj_204 (.A(cnt_init[0]), .B(num1_delay[15]), .C(n25559), 
         .D(n25650), .Z(num1_delay_15__N_780[15])) /* synthesis lut_function=(A (B (D))+!A (B (C+(D)))) */ ;
    defparam i1_4_lut_adj_204.init = 16'hcc40;
    LUT4 cnt_main_0__bdd_4_lut_21655 (.A(cnt_main[1]), .B(cnt_main[2]), 
         .C(time_data[20]), .D(time_data[8]), .Z(n24695)) /* synthesis lut_function=(!(A+!(B (D)+!B (C)))) */ ;
    defparam cnt_main_0__bdd_4_lut_21655.init = 16'h5410;
    LUT4 i2_4_lut_adj_205 (.A(n9753), .B(state[2]), .C(n35), .D(n31_adj_5153), 
         .Z(state_back_5__N_659[1])) /* synthesis lut_function=(A+(B (C)+!B (C+(D)))) */ ;
    defparam i2_4_lut_adj_205.init = 16'hfbfa;
    LUT4 i1_4_lut_adj_206 (.A(state[0]), .B(n16443), .C(state[2]), .D(state_back_5__N_858[1]), 
         .Z(n9753)) /* synthesis lut_function=(!(A (B+(C))+!A (B+!(C (D))))) */ ;
    defparam i1_4_lut_adj_206.init = 16'h1202;
    LUT4 i1_4_lut_adj_207 (.A(state_back[1]), .B(state[0]), .C(n25653), 
         .D(n24_adj_5154), .Z(n35)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_207.init = 16'haaa8;
    LUT4 i50_4_lut (.A(state_back[1]), .B(n25586), .C(state[3]), .D(n25649), 
         .Z(n31_adj_5153)) /* synthesis lut_function=(!((B (C)+!B (C (D)))+!A)) */ ;
    defparam i50_4_lut.init = 16'h0a2a;
    LUT4 i1_4_lut_adj_208 (.A(cnt_init[0]), .B(state_back[1]), .C(n25559), 
         .D(n25650), .Z(state_back_5__N_858[1])) /* synthesis lut_function=(A (B (D))+!A (B (C+(D)))) */ ;
    defparam i1_4_lut_adj_208.init = 16'hcc40;
    LUT4 i1_2_lut_adj_209 (.A(state[3]), .B(state[2]), .Z(n24_adj_5154)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_209.init = 16'h8888;
    LUT4 i73_2_lut_rep_409 (.A(state[2]), .B(state[3]), .Z(n25691)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i73_2_lut_rep_409.init = 16'h6666;
    LUT4 i1_2_lut_rep_311_3_lut_4_lut_4_lut (.A(state[2]), .B(state[3]), 
         .C(n25695), .D(n25760), .Z(n25593)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_2_lut_rep_311_3_lut_4_lut_4_lut.init = 16'h0004;
    LUT4 i1_3_lut_rep_354_4_lut (.A(state[2]), .B(state[3]), .C(n25754), 
         .D(n42_adj_5155), .Z(n25636)) /* synthesis lut_function=(A (B (D)+!B ((D)+!C))+!A (B ((D)+!C)+!B (D))) */ ;
    defparam i1_3_lut_rep_354_4_lut.init = 16'hff06;
    LUT4 i1_4_lut_adj_210 (.A(n24_adj_5156), .B(state_back[2]), .C(n25649), 
         .D(n9_adj_5058), .Z(state_back_5__N_659[2])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A ((D)+!B))) */ ;
    defparam i1_4_lut_adj_210.init = 16'h0ace;
    LUT4 i1_2_lut_rep_327_3_lut_4_lut (.A(state[2]), .B(state[3]), .C(n25695), 
         .D(n25760), .Z(n25609)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A ((C+(D))+!B))) */ ;
    defparam i1_2_lut_rep_327_3_lut_4_lut.init = 16'h0006;
    LUT4 i1_4_lut_adj_211 (.A(n25326), .B(state_back[3]), .C(n25649), 
         .D(n9_adj_5058), .Z(state_back_5__N_659[3])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A ((D)+!B))) */ ;
    defparam i1_4_lut_adj_211.init = 16'h0ace;
    LUT4 i1_4_lut_adj_212 (.A(n24_adj_5157), .B(state_back[4]), .C(n25649), 
         .D(n9_adj_5058), .Z(state_back_5__N_659[4])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A ((D)+!B))) */ ;
    defparam i1_4_lut_adj_212.init = 16'h0ace;
    LUT4 i1_4_lut_adj_213 (.A(n24_adj_5158), .B(state_back[5]), .C(n25649), 
         .D(n9_adj_5058), .Z(state_back_5__N_659[5])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A ((D)+!B))) */ ;
    defparam i1_4_lut_adj_213.init = 16'h0ace;
    LUT4 i2_2_lut_3_lut_4_lut_4_lut (.A(state[2]), .B(state[3]), .C(cnt_scan[3]), 
         .D(n25649), .Z(n6_adj_5101)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i2_2_lut_3_lut_4_lut_4_lut.init = 16'h0040;
    LUT4 i20789_2_lut_rep_410 (.A(state[1]), .B(state[5]), .Z(n25692)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i20789_2_lut_rep_410.init = 16'heeee;
    LUT4 i13252_4_lut_4_lut (.A(num1[0]), .B(n1359), .C(n1358), .D(n1357), 
         .Z(n93)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C (D)))+!A ((C+!(D))+!B))) */ ;
    defparam i13252_4_lut_4_lut.init = 16'h2c00;
    LUT4 i20911_2_lut_3_lut (.A(state[1]), .B(state[5]), .C(n23674), .Z(n23787)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i20911_2_lut_3_lut.init = 16'hfefe;
    LUT4 i13072_2_lut_rep_411 (.A(state[3]), .B(state[2]), .Z(n25693)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i13072_2_lut_rep_411.init = 16'heeee;
    LUT4 cnt_main_0__bdd_4_lut_21749 (.A(cnt_main[1]), .B(cnt_main[2]), 
         .C(time_data[16]), .D(time_data[12]), .Z(n24696)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)))) */ ;
    defparam cnt_main_0__bdd_4_lut_21749.init = 16'h6420;
    LUT4 i2_3_lut_4_lut_adj_214 (.A(state[3]), .B(state[2]), .C(state[4]), 
         .D(state[0]), .Z(n42_adj_5155)) /* synthesis lut_function=(!(A+(B+(C (D)+!C !(D))))) */ ;
    defparam i2_3_lut_4_lut_adj_214.init = 16'h0110;
    LUT4 i1_4_lut_adj_215 (.A(n25585), .B(n14556), .C(n29), .D(state[3]), 
         .Z(clk_c_enable_1432)) /* synthesis lut_function=(A (B)+!A (B+(C (D)))) */ ;
    defparam i1_4_lut_adj_215.init = 16'hdccc;
    LUT4 i2_4_lut_adj_216 (.A(n29), .B(num1_7__N_724[3]), .C(state[3]), 
         .D(state[0]), .Z(n14556)) /* synthesis lut_function=(!((B (C)+!B (C+!(D)))+!A)) */ ;
    defparam i2_4_lut_adj_216.init = 16'h0a08;
    LUT4 i1878_2_lut (.A(state[1]), .B(state[0]), .Z(n10049)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1878_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_rep_412 (.A(cnt_write[3]), .B(cnt_write[2]), .Z(n25694)) /* synthesis lut_function=(A+(B)) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(147[7] 167[14])
    defparam i1_2_lut_rep_412.init = 16'heeee;
    LUT4 i21448_4_lut (.A(state[0]), .B(n19_adj_5092), .C(n24_adj_5159), 
         .D(x_ph[1]), .Z(x_ph_7__N_519[1])) /* synthesis lut_function=(A ((D)+!B)+!A !(B (C+!(D))+!B (C))) */ ;
    defparam i21448_4_lut.init = 16'haf23;
    LUT4 i15039_4_lut (.A(x_ph[1]), .B(n89), .C(state[1]), .D(n94), 
         .Z(n24_adj_5159)) /* synthesis lut_function=(A (B (C (D)))+!A (B+!(C))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(29[13:18])
    defparam i15039_4_lut.init = 16'hc545;
    LUT4 i1_2_lut_rep_400_3_lut (.A(cnt_write[3]), .B(cnt_write[2]), .C(cnt_write[1]), 
         .Z(n25682)) /* synthesis lut_function=(A+(B+(C))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(147[7] 167[14])
    defparam i1_2_lut_rep_400_3_lut.init = 16'hfefe;
    LUT4 i1_3_lut_adj_217 (.A(n20788), .B(n83), .C(x_ph[2]), .Z(x_ph_7__N_519[2])) /* synthesis lut_function=(!(A (B)+!A !((C)+!B))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(29[13:18])
    defparam i1_3_lut_adj_217.init = 16'h7373;
    LUT4 i66_4_lut_4_lut (.A(cnt_main[1]), .B(time_data[11]), .C(cnt_main[2]), 
         .D(time_data[23]), .Z(n45)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(58[8:12])
    defparam i66_4_lut_4_lut.init = 16'h4f40;
    LUT4 i13137_2_lut_rep_413 (.A(state[1]), .B(state[0]), .Z(n25695)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i13137_2_lut_rep_413.init = 16'heeee;
    LUT4 n23706_bdd_2_lut_3_lut_4_lut_4_lut_4_lut (.A(n25676), .B(n25753), 
         .C(n25601), .D(n25635), .Z(n25119)) /* synthesis lut_function=(A (C+!(D))+!A (B (C)+!B (C+!(D)))) */ ;
    defparam n23706_bdd_2_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hf0fb;
    LUT4 i13877_2_lut_3_lut_4_lut (.A(state[1]), .B(state[0]), .C(n2557), 
         .D(n25605), .Z(n16664)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D)))) */ ;
    defparam i13877_2_lut_3_lut_4_lut.init = 16'heee0;
    LUT4 cnt_scan_2__bdd_3_lut_22024 (.A(x_pl[4]), .B(cnt_scan[0]), .C(cnt_scan[1]), 
         .Z(n24711)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam cnt_scan_2__bdd_3_lut_22024.init = 16'h8080;
    LUT4 i21442_4_lut (.A(state[0]), .B(x_ph[3]), .C(n24_adj_5160), .D(n19_adj_5092), 
         .Z(x_ph_7__N_519[3])) /* synthesis lut_function=(A (B+!(D))+!A !(B (C)+!B (C+(D)))) */ ;
    defparam i21442_4_lut.init = 16'h8caf;
    LUT4 i41_4_lut_adj_218 (.A(x_ph[3]), .B(n23318), .C(state[1]), .D(n4_adj_5161), 
         .Z(n24_adj_5160)) /* synthesis lut_function=(A (B (C (D)))+!A (B ((D)+!C)+!B !(C))) */ ;
    defparam i41_4_lut_adj_218.init = 16'hc505;
    LUT4 i21477_2_lut_rep_414 (.A(state[2]), .B(state[0]), .Z(n25696)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i21477_2_lut_rep_414.init = 16'h1111;
    LUT4 i2_3_lut_rep_353 (.A(num2[3]), .B(char[3]), .C(n6_adj_5088), 
         .Z(n25635)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B (C)+!B !(C)))) */ ;
    defparam i2_3_lut_rep_353.init = 16'h6969;
    LUT4 i1_2_lut_rep_415 (.A(cnt_init[2]), .B(cnt_init[1]), .Z(n25697)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut_rep_415.init = 16'h2222;
    LUT4 cnt_scan_2__bdd_3_lut_21664 (.A(x_ph[4]), .B(cnt_scan[0]), .C(cnt_scan[1]), 
         .Z(n24710)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;
    defparam cnt_scan_2__bdd_3_lut_21664.init = 16'h0202;
    LUT4 i1_2_lut_rep_288_3_lut_4_lut (.A(cnt_init[2]), .B(cnt_init[1]), 
         .C(oled_dcn_N_888), .D(n25698), .Z(n25570)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_rep_288_3_lut_4_lut.init = 16'h0020;
    LUT4 i21432_4_lut (.A(state[0]), .B(x_ph[4]), .C(n24_adj_5162), .D(n19_adj_5092), 
         .Z(x_ph_7__N_519[4])) /* synthesis lut_function=(A (B+!(D))+!A !(B (C)+!B (C+(D)))) */ ;
    defparam i21432_4_lut.init = 16'h8caf;
    LUT4 i41_4_lut_adj_219 (.A(x_ph[4]), .B(n9), .C(state[1]), .D(n4_adj_5057), 
         .Z(n24_adj_5162)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A !((D)+!C))) */ ;
    defparam i41_4_lut_adj_219.init = 16'h7505;
    LUT4 n3_bdd_3_lut_21705 (.A(cnt_main[2]), .B(cnt_main[1]), .C(\tamp_data[6] ), 
         .Z(n24714)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam n3_bdd_3_lut_21705.init = 16'h8080;
    LUT4 i21429_4_lut (.A(state[0]), .B(x_ph[5]), .C(n24_adj_5163), .D(n19_adj_5092), 
         .Z(x_ph_7__N_519[5])) /* synthesis lut_function=(A (B+!(D))+!A !(B (C)+!B (C+(D)))) */ ;
    defparam i21429_4_lut.init = 16'h8caf;
    LUT4 i41_4_lut_adj_220 (.A(x_ph[5]), .B(n23318), .C(state[1]), .D(n4_adj_5078), 
         .Z(n24_adj_5163)) /* synthesis lut_function=(A (B (C (D)))+!A (B ((D)+!C)+!B !(C))) */ ;
    defparam i41_4_lut_adj_220.init = 16'hc505;
    LUT4 i1_2_lut_3_lut_adj_221 (.A(cnt_init[2]), .B(cnt_init[1]), .C(cnt_init[0]), 
         .Z(n4_adj_5115)) /* synthesis lut_function=(A ((C)+!B)+!A (C)) */ ;
    defparam i1_2_lut_3_lut_adj_221.init = 16'hf2f2;
    LUT4 i1_3_lut_adj_222 (.A(n20788), .B(n83), .C(x_ph[6]), .Z(x_ph_7__N_519[6])) /* synthesis lut_function=(!(A (B)+!A !((C)+!B))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(29[13:18])
    defparam i1_3_lut_adj_222.init = 16'h7373;
    LUT4 i13163_2_lut_rep_416 (.A(cnt_init[4]), .B(cnt_init[3]), .Z(n25698)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i13163_2_lut_rep_416.init = 16'heeee;
    LUT4 i1_2_lut_rep_369_3_lut_4_lut (.A(cnt_init[4]), .B(cnt_init[3]), 
         .C(cnt_init[1]), .D(cnt_init[2]), .Z(n25651)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_2_lut_rep_369_3_lut_4_lut.init = 16'h0100;
    LUT4 i7_4_lut_adj_223 (.A(num2[0]), .B(n14_adj_5164), .C(n10_adj_5165), 
         .D(num2[6]), .Z(n322)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(106[11:15])
    defparam i7_4_lut_adj_223.init = 16'hfffe;
    LUT4 i1_2_lut_rep_383_3_lut (.A(cnt_init[4]), .B(cnt_init[3]), .C(state[2]), 
         .Z(n25665)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_rep_383_3_lut.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_4_lut_adj_224 (.A(cnt_init[4]), .B(cnt_init[3]), 
         .C(n23755), .D(state[2]), .Z(n4434)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_224.init = 16'h0100;
    LUT4 i6_4_lut_adj_225 (.A(num2[3]), .B(num2[1]), .C(num2[5]), .D(num2[7]), 
         .Z(n14_adj_5164)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(106[11:15])
    defparam i6_4_lut_adj_225.init = 16'hfffe;
    LUT4 i1_2_lut_4_lut_adj_226 (.A(num2[3]), .B(char[3]), .C(n6_adj_5088), 
         .D(num2[0]), .Z(n4_adj_5148)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C+(D)))+!A (B (C+(D))+!B ((D)+!C))) */ ;
    defparam i1_2_lut_4_lut_adj_226.init = 16'hff69;
    LUT4 i1_2_lut_3_lut_adj_227 (.A(cnt_scan[0]), .B(cnt_scan[1]), .C(x_ph[2]), 
         .Z(n4_adj_5087)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(111[7] 142[14])
    defparam i1_2_lut_3_lut_adj_227.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_228 (.A(cnt_scan[0]), .B(cnt_scan[1]), .C(x_ph[6]), 
         .Z(n69)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(111[7] 142[14])
    defparam i1_2_lut_3_lut_adj_228.init = 16'h1010;
    LUT4 i2_2_lut_adj_229 (.A(num2[2]), .B(num2[4]), .Z(n10_adj_5165)) /* synthesis lut_function=(A+(B)) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(106[11:15])
    defparam i2_2_lut_adj_229.init = 16'heeee;
    LUT4 n26041_bdd_2_lut (.A(n26777), .B(state[1]), .Z(n26042)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam n26041_bdd_2_lut.init = 16'h2222;
    LUT4 n25060_bdd_3_lut_21938 (.A(n8855), .B(cnt_scan[0]), .C(num2[0]), 
         .Z(n25211)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;
    defparam n25060_bdd_3_lut_21938.init = 16'h0101;
    LUT4 i13538_2_lut (.A(x_ph[1]), .B(cnt_scan[0]), .Z(n4)) /* synthesis lut_function=(A+(B)) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(111[7] 142[14])
    defparam i13538_2_lut.init = 16'heeee;
    CCU2D add_143_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt_delay[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n20497), .S1(n2559[0]));   // g:/fpga/mxo2/system/project/oled12832.v(172[29:45])
    defparam add_143_1.INIT0 = 16'hF000;
    defparam add_143_1.INIT1 = 16'h5555;
    defparam add_143_1.INJECT1_0 = "NO";
    defparam add_143_1.INJECT1_1 = "NO";
    LUT4 n25060_bdd_2_lut (.A(n25060), .B(n1354), .Z(n25212)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam n25060_bdd_2_lut.init = 16'h2222;
    LUT4 i1_3_lut_4_lut_adj_230 (.A(n25711), .B(n25763), .C(n9), .D(x_ph[3]), 
         .Z(n4_adj_5161)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A (C (D)))) */ ;
    defparam i1_3_lut_4_lut_adj_230.init = 16'h0ddd;
    LUT4 n25060_bdd_3_lut (.A(n25063), .B(n25064), .C(n1354), .Z(n25213)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n25060_bdd_3_lut.init = 16'hacac;
    LUT4 i1_2_lut_rep_363_2_lut (.A(cnt_main[4]), .B(cnt_main[2]), .Z(n25645)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut_rep_363_2_lut.init = 16'h4444;
    LUT4 i2_4_lut_4_lut (.A(cnt_main[4]), .B(time_data[2]), .C(cnt_main[1]), 
         .D(cnt_main[3]), .Z(n20744)) /* synthesis lut_function=(!(A+!(B (D)+!B (C (D))))) */ ;
    defparam i2_4_lut_4_lut.init = 16'h5400;
    LUT4 i1_2_lut_rep_297 (.A(n1354), .B(n1356), .Z(n25579)) /* synthesis lut_function=(A (B)) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(129[51:75])
    defparam i1_2_lut_rep_297.init = 16'h8888;
    LUT4 i1_4_lut_4_lut_adj_231 (.A(cnt_main[4]), .B(n68_adj_5114), .C(n25631), 
         .D(char[3]), .Z(n4_adj_5113)) /* synthesis lut_function=(A (C (D))+!A (B+(C (D)))) */ ;
    defparam i1_4_lut_4_lut_adj_231.init = 16'hf444;
    LUT4 i1_4_lut_4_lut_adj_232 (.A(cnt_main[4]), .B(cnt_main[1]), .C(n99), 
         .D(n105), .Z(n89_adj_5118)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;
    defparam i1_4_lut_4_lut_adj_232.init = 16'h5140;
    LUT4 i1_4_lut_4_lut_adj_233 (.A(cnt_main[4]), .B(n25762), .C(n39), 
         .D(n25786), .Z(n4_adj_5107)) /* synthesis lut_function=(A (B (D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_4_lut_adj_233.init = 16'hdc50;
    LUT4 i1_4_lut_4_lut_adj_234 (.A(cnt_main[4]), .B(n43), .C(n41_adj_5109), 
         .D(n16111), .Z(char_7__N_756[2])) /* synthesis lut_function=(A (C+!(D))+!A (B+(C+!(D)))) */ ;
    defparam i1_4_lut_4_lut_adj_234.init = 16'hf4ff;
    LUT4 i110_2_lut_2_lut (.A(cnt_main[4]), .B(n58), .Z(n94)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i110_2_lut_2_lut.init = 16'h4444;
    PFUMX i21028 (.BLUT(n23903), .ALUT(n23904), .C0(cnt_scan[4]), .Z(char_reg_7__N_772[5]));
    LUT4 i20671_2_lut_rep_312_4_lut (.A(num2[3]), .B(char[3]), .C(n6_adj_5088), 
         .D(n25676), .Z(n25594)) /* synthesis lut_function=(A (B (C (D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C (D)))) */ ;
    defparam i20671_2_lut_rep_312_4_lut.init = 16'h9600;
    LUT4 i1_2_lut_3_lut_adj_235 (.A(cnt_main[1]), .B(cnt_main[3]), .C(char[3]), 
         .Z(n9872)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_235.init = 16'h1010;
    PFUMX i21802 (.BLUT(n24963), .ALUT(n24962), .C0(n25635), .Z(n24964));
    PFUMX i21016 (.BLUT(n23891), .ALUT(n23892), .C0(cnt_scan[4]), .Z(char_reg_7__N_772[3]));
    LUT4 i13529_3_lut (.A(x_ph[5]), .B(cnt_scan[1]), .C(cnt_scan[0]), 
         .Z(n6_adj_5059)) /* synthesis lut_function=(!(A (B)+!A (B+!(C)))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(111[7] 142[14])
    defparam i13529_3_lut.init = 16'h3232;
    LUT4 mux_131_Mux_1_i11_3_lut_4_lut (.A(num1[0]), .B(n25557), .C(cnt_scan[0]), 
         .D(n864), .Z(n11_adj_5166)) /* synthesis lut_function=(!(A (C+!(D))+!A (B (C+!(D))+!B !(C+(D))))) */ ;
    defparam mux_131_Mux_1_i11_3_lut_4_lut.init = 16'h1f10;
    LUT4 i1_2_lut_4_lut_adj_236 (.A(n25691), .B(n42_adj_5155), .C(n25754), 
         .D(n25692), .Z(n20715)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A ((D)+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_236.init = 16'h00ce;
    LUT4 n26039_bdd_4_lut (.A(n26039), .B(n27), .C(state[3]), .D(state[0]), 
         .Z(n26777)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam n26039_bdd_4_lut.init = 16'h00ca;
    PFUMX i21019 (.BLUT(n23894), .ALUT(n23895), .C0(cnt_scan[4]), .Z(char_reg_7__N_772[2]));
    FD1P3AX oled_dat_372 (.D(n20727), .SP(clk_c_enable_1421), .CK(clk_c), 
            .Q(oled_dat_c)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam oled_dat_372.GSR = "ENABLED";
    LUT4 mux_1250_i1_4_lut (.A(n30_adj_5167), .B(char_reg_7__N_772[0]), 
         .C(state[3]), .D(n23821), .Z(n3492[0])) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B ((D)+!C))) */ ;
    defparam mux_1250_i1_4_lut.init = 16'hccac;
    PFUMX i21031 (.BLUT(n23906), .ALUT(n23907), .C0(cnt_scan[4]), .Z(char_reg_7__N_772[4]));
    PFUMX i22165 (.BLUT(n25787), .ALUT(n25788), .C0(state[0]), .Z(n25789));
    LUT4 mux_131_Mux_0_i31_4_lut (.A(n18_adj_5168), .B(n25826), .C(state[3]), 
         .D(n25558), .Z(char_reg_7__N_772[0])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A !((C+!(D))+!B)) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(111[7] 142[14])
    defparam mux_131_Mux_0_i31_4_lut.init = 16'haca0;
    LUT4 cnt_write_4__bdd_3_lut_21903_4_lut (.A(cnt_write[0]), .B(n25682), 
         .C(state[4]), .D(cnt_write[4]), .Z(n25115)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C (D))))) */ ;
    defparam cnt_write_4__bdd_3_lut_21903_4_lut.init = 16'h10e0;
    FD1P3AY oled_clk_371 (.D(n22465), .SP(clk_c_enable_1423), .CK(clk_c), 
            .Q(oled_clk_c)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam oled_clk_371.GSR = "ENABLED";
    LUT4 i21473_4_lut (.A(n50), .B(n24187), .C(n25693), .D(n25695), 
         .Z(n42)) /* synthesis lut_function=(A (B (C+(D)))+!A (B)) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(41[4] 175[11])
    defparam i21473_4_lut.init = 16'hccc4;
    LUT4 i21472_4_lut (.A(n44), .B(n25760), .C(n26042), .D(n25693), 
         .Z(n24187)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B+!(C))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(41[4] 175[11])
    defparam i21472_4_lut.init = 16'hcfcd;
    LUT4 i72_4_lut (.A(state[0]), .B(n36), .C(state[1]), .D(n25610), 
         .Z(n44)) /* synthesis lut_function=(!(A (C)+!A (B ((D)+!C)+!B !(C)))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(41[4] 175[11])
    defparam i72_4_lut.init = 16'h1a5a;
    PFUMX i21022 (.BLUT(n23897), .ALUT(n23898), .C0(cnt_scan[4]), .Z(char_reg_7__N_772[1]));
    LUT4 i20944_3_lut (.A(cnt_scan[4]), .B(cnt_scan[3]), .C(cnt_scan[2]), 
         .Z(n23821)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(111[7] 142[14])
    defparam i20944_3_lut.init = 16'h0202;
    LUT4 i3_3_lut_rep_284_4_lut (.A(n1354), .B(n1356), .C(n1357), .D(n1355), 
         .Z(n25566)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(129[51:75])
    defparam i3_3_lut_rep_284_4_lut.init = 16'h0080;
    L6MUX21 i21051 (.D0(n23953), .D1(n20_adj_5169), .SD(cnt_scan[1]), 
            .Z(n23928));
    LUT4 n2533_bdd_4_lut_4_lut (.A(cnt_write[0]), .B(n25682), .C(cnt_write[4]), 
         .D(state[4]), .Z(n25496)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam n2533_bdd_4_lut_4_lut.init = 16'h2000;
    L6MUX21 mux_131_Mux_0_i30 (.D0(n22_adj_5170), .D1(n23935), .SD(n25748), 
            .Z(n30_adj_5167)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;
    PFUMX mux_131_Mux_5_i20 (.BLUT(n6170), .ALUT(n2162[21]), .C0(n23867), 
          .Z(n20_adj_5169)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;
    CCU2D add_2997_7 (.A0(char[5]), .B0(n25671), .C0(num1[5]), .D0(GND_net), 
          .A1(char[6]), .B1(n23153), .C1(num1[6]), .D1(GND_net), .CIN(n20573), 
          .S0(n1355), .S1(n1354));   // g:/fpga/mxo2/system/project/oled12832.v(129[56:62])
    defparam add_2997_7.INIT0 = 16'h9969;
    defparam add_2997_7.INIT1 = 16'h9969;
    defparam add_2997_7.INJECT1_0 = "NO";
    defparam add_2997_7.INJECT1_1 = "NO";
    CCU2D add_2997_5 (.A0(char[3]), .B0(n25745), .C0(num1[3]), .D0(GND_net), 
          .A1(char[4]), .B1(n20442), .C1(num1[4]), .D1(GND_net), .CIN(n20572), 
          .COUT(n20573), .S0(n1357), .S1(n1356));   // g:/fpga/mxo2/system/project/oled12832.v(129[56:62])
    defparam add_2997_5.INIT0 = 16'h9969;
    defparam add_2997_5.INIT1 = 16'h9969;
    defparam add_2997_5.INJECT1_0 = "NO";
    defparam add_2997_5.INJECT1_1 = "NO";
    LUT4 i21599_2_lut_3_lut_4_lut_1_lut (.A(cnt_main[0]), .Z(n2[0])) /* synthesis lut_function=(!(A)) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(58[8:12])
    defparam i21599_2_lut_3_lut_4_lut_1_lut.init = 16'h5555;
    LUT4 i2_3_lut_4_lut_adj_237 (.A(n1354), .B(n1356), .C(n1355), .D(n1357), 
         .Z(n23134)) /* synthesis lut_function=(((C+!(D))+!B)+!A) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(129[51:75])
    defparam i2_3_lut_4_lut_adj_237.init = 16'hf7ff;
    CCU2D add_38_17 (.A0(cnt_c[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n20496), 
          .S0(n141[15]));   // g:/fpga/mxo2/system/project/oled12832.v(88[19:29])
    defparam add_38_17.INIT0 = 16'h5aaa;
    defparam add_38_17.INIT1 = 16'h0000;
    defparam add_38_17.INJECT1_0 = "NO";
    defparam add_38_17.INJECT1_1 = "NO";
    LUT4 i1_4_lut_4_lut_adj_238 (.A(cnt_main[0]), .B(cnt_main[1]), .C(n25763), 
         .D(n25798), .Z(n4_adj_5096)) /* synthesis lut_function=(!(A+!(B ((D)+!C)+!B (D)))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(58[8:12])
    defparam i1_4_lut_4_lut_adj_238.init = 16'h5504;
    LUT4 i1_2_lut_rep_429 (.A(cnt_main[1]), .B(cnt_main[0]), .Z(n25711)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_429.init = 16'h8888;
    LUT4 i1_3_lut_4_lut_adj_239 (.A(cnt_main[1]), .B(cnt_main[0]), .C(n25743), 
         .D(cnt_main[4]), .Z(n36)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;
    defparam i1_3_lut_4_lut_adj_239.init = 16'hff80;
    LUT4 i2_3_lut_rep_322_4_lut (.A(state[3]), .B(n25683), .C(state[5]), 
         .D(state[4]), .Z(n25604)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(169[5:10])
    defparam i2_3_lut_rep_322_4_lut.init = 16'hfeff;
    LUT4 i1_4_lut_3_lut (.A(cnt_main[1]), .B(n25629), .C(n25718), .Z(n16632)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i1_4_lut_3_lut.init = 16'he4e4;
    LUT4 i13076_2_lut_rep_431 (.A(state[3]), .B(state[0]), .Z(n25713)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i13076_2_lut_rep_431.init = 16'heeee;
    LUT4 i30_4_lut_3_lut (.A(state[3]), .B(state[0]), .C(state[1]), .Z(n17_adj_5171)) /* synthesis lut_function=(!(A (B+(C))+!A (B (C)+!B !(C)))) */ ;
    defparam i30_4_lut_3_lut.init = 16'h1616;
    LUT4 i13613_2_lut_3_lut (.A(state[3]), .B(state[0]), .C(num1_7__N_724[3]), 
         .Z(n16391)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i13613_2_lut_3_lut.init = 16'hfefe;
    LUT4 i21467_4_lut (.A(state[0]), .B(num1_delay[0]), .C(n24_adj_5172), 
         .D(n27_adj_5133), .Z(num1_delay_15__N_605[0])) /* synthesis lut_function=(A (B+!(D))+!A !(B (C)+!B (C+(D)))) */ ;
    defparam i21467_4_lut.init = 16'h8caf;
    LUT4 i2_3_lut_rep_323_4_lut (.A(state[3]), .B(n25683), .C(state[5]), 
         .D(state[4]), .Z(n25605)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(169[5:10])
    defparam i2_3_lut_rep_323_4_lut.init = 16'hffef;
    CCU2D add_2997_3 (.A0(char[1]), .B0(num1[1]), .C0(GND_net), .D0(GND_net), 
          .A1(char[1]), .B1(char[2]), .C1(num1[2]), .D1(GND_net), .CIN(n20571), 
          .COUT(n20572), .S0(n1359), .S1(n1358));   // g:/fpga/mxo2/system/project/oled12832.v(129[56:62])
    defparam add_2997_3.INIT0 = 16'ha666;
    defparam add_2997_3.INIT1 = 16'h6696;
    defparam add_2997_3.INJECT1_0 = "NO";
    defparam add_2997_3.INJECT1_1 = "NO";
    LUT4 i21865_then_4_lut (.A(cnt_main[2]), .B(cnt_main[4]), .C(cnt_main[1]), 
         .D(cnt_main[3]), .Z(n25797)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A (B (C+(D))+!B (D)))) */ ;
    defparam i21865_then_4_lut.init = 16'h201f;
    CCU2D add_38_15 (.A0(cnt_c[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt_c[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n20495), .COUT(n20496), .S0(n141[13]), .S1(n141[14]));   // g:/fpga/mxo2/system/project/oled12832.v(88[19:29])
    defparam add_38_15.INIT0 = 16'h5aaa;
    defparam add_38_15.INIT1 = 16'h5aaa;
    defparam add_38_15.INJECT1_0 = "NO";
    defparam add_38_15.INJECT1_1 = "NO";
    FD1P3AX oled_dcn_370 (.D(n23342), .SP(clk_c_enable_1427), .CK(clk_c), 
            .Q(oled_dcn_c)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam oled_dcn_370.GSR = "ENABLED";
    LUT4 i21865_else_4_lut (.A(cnt_main[2]), .B(cnt_main[4]), .C(cnt_main[1]), 
         .D(cnt_main[3]), .Z(n25796)) /* synthesis lut_function=(!(A (B+!(C (D)+!C !(D)))+!A (B+((D)+!C)))) */ ;
    defparam i21865_else_4_lut.init = 16'h2012;
    LUT4 i2_3_lut_rep_436 (.A(cnt_main[3]), .B(cnt_main[4]), .C(cnt_main[2]), 
         .Z(n25718)) /* synthesis lut_function=((B+(C))+!A) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(65[8:12])
    defparam i2_3_lut_rep_436.init = 16'hfdfd;
    LUT4 i2_3_lut_3_lut_4_lut (.A(cnt_scan[1]), .B(cnt_scan[0]), .C(cnt_scan[4]), 
         .D(cnt_scan[2]), .Z(n20791)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (((D)+!C)+!B))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(110[42:57])
    defparam i2_3_lut_3_lut_4_lut.init = 16'h0060;
    LUT4 mux_1283_i2_3_lut_4_lut (.A(cnt_scan[1]), .B(cnt_scan[0]), .C(n3599), 
         .D(n4264[1]), .Z(cnt_scan_4__N_682[1])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(110[42:57])
    defparam mux_1283_i2_3_lut_4_lut.init = 16'hf606;
    LUT4 i13185_2_lut_rep_437 (.A(cnt_scan[0]), .B(cnt_scan[1]), .Z(n25719)) /* synthesis lut_function=(A (B)) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(111[7] 142[14])
    defparam i13185_2_lut_rep_437.init = 16'h8888;
    CCU2D add_2997_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(num1[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n20571));   // g:/fpga/mxo2/system/project/oled12832.v(129[56:62])
    defparam add_2997_1.INIT0 = 16'h0000;
    defparam add_2997_1.INIT1 = 16'h0aaa;
    defparam add_2997_1.INJECT1_0 = "NO";
    defparam add_2997_1.INJECT1_1 = "NO";
    PFUMX mux_131_Mux_0_i22 (.BLUT(n6550), .ALUT(n23349), .C0(cnt_scan[3]), 
          .Z(n22_adj_5170)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;
    LUT4 i2694_2_lut_3_lut_4_lut (.A(cnt_scan[0]), .B(cnt_scan[1]), .C(cnt_scan[3]), 
         .D(cnt_scan[2]), .Z(n331[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(111[7] 142[14])
    defparam i2694_2_lut_3_lut_4_lut.init = 16'h78f0;
    LUT4 i41_4_lut_adj_240 (.A(num1_delay[0]), .B(n16443), .C(state[2]), 
         .D(n23253), .Z(n24_adj_5172)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C)+!B !((D)+!C)))) */ ;
    defparam i41_4_lut_adj_240.init = 16'h3505;
    LUT4 i1_2_lut_3_lut_adj_241 (.A(cnt_scan[0]), .B(cnt_scan[1]), .C(x_pl[6]), 
         .Z(n68)) /* synthesis lut_function=(A (B (C))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(111[7] 142[14])
    defparam i1_2_lut_3_lut_adj_241.init = 16'h8080;
    PFUMX i47 (.BLUT(n6_adj_5075), .ALUT(n23280), .C0(state[3]), .Z(n24_adj_5156));
    LUT4 i94_4_lut_3_lut (.A(state[2]), .B(state[0]), .C(n25581), .Z(n69_adj_5173)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(41[4] 175[11])
    defparam i94_4_lut_3_lut.init = 16'h6464;
    L6MUX21 i29 (.D0(n13_adj_5174), .D1(n23947), .SD(cnt_scan[2]), .Z(n16_adj_5130));
    LUT4 i1_4_lut_adj_242 (.A(cnt_write[1]), .B(cnt_write[4]), .C(cnt_write[0]), 
         .D(n25694), .Z(n23223)) /* synthesis lut_function=(!(A+(B ((D)+!C)+!B (C+(D))))) */ ;
    defparam i1_4_lut_adj_242.init = 16'h0041;
    LUT4 i13092_2_lut_rep_478 (.A(state[5]), .B(state[4]), .Z(n25760)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i13092_2_lut_rep_478.init = 16'heeee;
    PFUMX i21768 (.BLUT(n24906), .ALUT(n24905), .C0(n1357), .Z(n24907));
    LUT4 i21493_2_lut_rep_276_4_lut (.A(n25678), .B(oled_dcn_N_888), .C(cnt_init[0]), 
         .D(state[0]), .Z(n25558)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i21493_2_lut_rep_276_4_lut.init = 16'h0001;
    LUT4 i1_2_lut_2_lut_adj_243 (.A(cnt_init[0]), .B(cnt_init[1]), .Z(n4_adj_5116)) /* synthesis lut_function=(!(A+!(B))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(79[49:64])
    defparam i1_2_lut_2_lut_adj_243.init = 16'h4444;
    LUT4 i1_2_lut_3_lut_4_lut_adj_244 (.A(n25760), .B(n25693), .C(n15856), 
         .D(n16743), .Z(n23318)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_244.init = 16'h1000;
    LUT4 i1_4_lut_4_lut_adj_245 (.A(n25678), .B(oled_dcn_N_888), .C(cnt_init[0]), 
         .D(n25677), .Z(n13)) /* synthesis lut_function=(A (D)+!A !(B+(C))) */ ;
    defparam i1_4_lut_4_lut_adj_245.init = 16'hab01;
    PFUMX mux_131_Mux_2_i18 (.BLUT(n16_adj_5136), .ALUT(n17_adj_5044), .C0(cnt_scan[1]), 
          .Z(n18_adj_5082)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;
    LUT4 n23548_bdd_4_lut_22003_4_lut (.A(cnt_init[0]), .B(state_back[3]), 
         .C(n25650), .D(n25559), .Z(n25324)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D)))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(79[49:64])
    defparam n23548_bdd_4_lut_22003_4_lut.init = 16'hc4c0;
    LUT4 i1_3_lut_rep_326_4_lut (.A(n25760), .B(n25693), .C(state[1]), 
         .D(state[0]), .Z(n25608)) /* synthesis lut_function=(!(A+(B+(C (D)+!C !(D))))) */ ;
    defparam i1_3_lut_rep_326_4_lut.init = 16'h0110;
    CCU2D add_38_13 (.A0(cnt_c[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt_c[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n20494), .COUT(n20495), .S0(n141[11]), .S1(n141[12]));   // g:/fpga/mxo2/system/project/oled12832.v(88[19:29])
    defparam add_38_13.INIT0 = 16'h5aaa;
    defparam add_38_13.INIT1 = 16'h5aaa;
    defparam add_38_13.INJECT1_0 = "NO";
    defparam add_38_13.INJECT1_1 = "NO";
    LUT4 i1772_2_lut_3_lut_4_lut (.A(n25760), .B(n25693), .C(state[1]), 
         .D(state[0]), .Z(n4432)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1772_2_lut_3_lut_4_lut.init = 16'h0100;
    CCU2D add_38_11 (.A0(cnt_c[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt_c[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n20493), .COUT(n20494), .S0(n141[9]), .S1(n141[10]));   // g:/fpga/mxo2/system/project/oled12832.v(88[19:29])
    defparam add_38_11.INIT0 = 16'h5aaa;
    defparam add_38_11.INIT1 = 16'h5aaa;
    defparam add_38_11.INJECT1_0 = "NO";
    defparam add_38_11.INJECT1_1 = "NO";
    LUT4 n2421_bdd_4_lut (.A(n23763), .B(n25601), .C(n25632), .D(n25635), 
         .Z(n25312)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C))+!A !(B (C+(D))+!B (C)))) */ ;
    defparam n2421_bdd_4_lut.init = 16'h74f0;
    CCU2D add_38_9 (.A0(cnt_c[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt_c[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n20492), 
          .COUT(n20493), .S0(n141[7]), .S1(n141[8]));   // g:/fpga/mxo2/system/project/oled12832.v(88[19:29])
    defparam add_38_9.INIT0 = 16'h5aaa;
    defparam add_38_9.INIT1 = 16'h5aaa;
    defparam add_38_9.INJECT1_0 = "NO";
    defparam add_38_9.INJECT1_1 = "NO";
    LUT4 i13593_2_lut_rep_367_3_lut_4_lut (.A(state[5]), .B(state[4]), .C(state[0]), 
         .D(state[1]), .Z(n25649)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13593_2_lut_rep_367_3_lut_4_lut.init = 16'hfffe;
    L6MUX21 i21034 (.D0(n23909), .D1(n23910), .SD(cnt_scan[2]), .Z(n23911));
    LUT4 mux_1090_i1_4_lut (.A(cnt_write[4]), .B(state[0]), .C(n25608), 
         .D(state[4]), .Z(n3153[0])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(41[4] 175[11])
    defparam mux_1090_i1_4_lut.init = 16'hcac0;
    L6MUX21 i21036 (.D0(n23956), .D1(n23959), .SD(cnt_scan[1]), .Z(n23913));
    L6MUX21 i21040 (.D0(n23915), .D1(n23916), .SD(cnt_scan[2]), .Z(n23917));
    L6MUX21 i21043 (.D0(n23918), .D1(n23919), .SD(cnt_scan[2]), .Z(n23920));
    LUT4 i1_2_lut_rep_274_4_lut (.A(n25579), .B(n1355), .C(n1357), .D(cnt_scan[0]), 
         .Z(n25556)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(129[51:75])
    defparam i1_2_lut_rep_274_4_lut.init = 16'h2000;
    LUT4 i1_4_lut_4_lut_adj_246 (.A(cnt_init[0]), .B(n23583), .C(n19_adj_5175), 
         .D(state[2]), .Z(n6_adj_5176)) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(79[49:64])
    defparam i1_4_lut_4_lut_adj_246.init = 16'hf400;
    LUT4 i2_4_lut_4_lut_4_lut (.A(cnt_init[0]), .B(state[4]), .C(n25677), 
         .D(n25651), .Z(n21246)) /* synthesis lut_function=(!(A+!(B ((D)+!C)))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(79[49:64])
    defparam i2_4_lut_4_lut_4_lut.init = 16'h4404;
    LUT4 i1_4_lut_4_lut_adj_247 (.A(cnt_init[0]), .B(n23581), .C(n19_adj_5177), 
         .D(state[2]), .Z(n6_adj_5178)) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(79[49:64])
    defparam i1_4_lut_4_lut_adj_247.init = 16'hf400;
    LUT4 i1_4_lut_then_4_lut (.A(cnt_main[4]), .B(cnt_main[2]), .C(cnt_main[3]), 
         .D(cnt_main[0]), .Z(n25801)) /* synthesis lut_function=(A+(B (C (D)))) */ ;
    defparam i1_4_lut_then_4_lut.init = 16'heaaa;
    CCU2D add_38_7 (.A0(cnt_c[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt_c[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n20491), 
          .COUT(n20492), .S0(n141[5]), .S1(n141[6]));   // g:/fpga/mxo2/system/project/oled12832.v(88[19:29])
    defparam add_38_7.INIT0 = 16'h5aaa;
    defparam add_38_7.INIT1 = 16'h5aaa;
    defparam add_38_7.INJECT1_0 = "NO";
    defparam add_38_7.INJECT1_1 = "NO";
    LUT4 i10770_4_lut_4_lut (.A(cnt_init[0]), .B(n25628), .C(n25651), 
         .D(state[4]), .Z(n13577)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A !(B (C+(D))+!B (C)))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(79[49:64])
    defparam i10770_4_lut_4_lut.init = 16'h5c50;
    L6MUX21 i21054 (.D0(n7110), .D1(n7112), .SD(cnt_scan[1]), .Z(n23931));
    LUT4 i1_4_lut_4_lut_adj_248 (.A(cnt_init[0]), .B(n25570), .C(n23312), 
         .D(n25628), .Z(n23314)) /* synthesis lut_function=(A (C (D))+!A (B (C)+!B (C (D)))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(79[49:64])
    defparam i1_4_lut_4_lut_adj_248.init = 16'hf040;
    LUT4 i1_4_lut_4_lut_adj_249 (.A(cnt_init[0]), .B(n23579), .C(n19_adj_5179), 
         .D(state[2]), .Z(n6_adj_5180)) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(79[49:64])
    defparam i1_4_lut_4_lut_adj_249.init = 16'hf400;
    LUT4 n2421_bdd_3_lut_22045 (.A(n23763), .B(n25601), .C(n25635), .Z(n25310)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam n2421_bdd_3_lut_22045.init = 16'h4040;
    LUT4 i2_3_lut_4_lut_adj_250 (.A(n25760), .B(n25693), .C(n16743), .D(n23157), 
         .Z(n89)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i2_3_lut_4_lut_adj_250.init = 16'h1000;
    LUT4 n25313_bdd_3_lut (.A(n25313), .B(n25310), .C(num2[0]), .Z(n25314)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25313_bdd_3_lut.init = 16'hcaca;
    CCU2D add_38_5 (.A0(cnt[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n20490), 
          .COUT(n20491), .S0(n141[3]), .S1(n141[4]));   // g:/fpga/mxo2/system/project/oled12832.v(88[19:29])
    defparam add_38_5.INIT0 = 16'h5aaa;
    defparam add_38_5.INIT1 = 16'h5aaa;
    defparam add_38_5.INJECT1_0 = "NO";
    defparam add_38_5.INJECT1_1 = "NO";
    CCU2D add_38_3 (.A0(cnt[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n20489), 
          .COUT(n20490), .S0(n141[1]), .S1(n141[2]));   // g:/fpga/mxo2/system/project/oled12832.v(88[19:29])
    defparam add_38_3.INIT0 = 16'h5aaa;
    defparam add_38_3.INIT1 = 16'h5aaa;
    defparam add_38_3.INJECT1_0 = "NO";
    defparam add_38_3.INJECT1_1 = "NO";
    CCU2D add_38_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n20489), 
          .S1(n141[0]));   // g:/fpga/mxo2/system/project/oled12832.v(88[19:29])
    defparam add_38_1.INIT0 = 16'hF000;
    defparam add_38_1.INIT1 = 16'h5555;
    defparam add_38_1.INJECT1_0 = "NO";
    defparam add_38_1.INJECT1_1 = "NO";
    LUT4 i1_4_lut_else_4_lut (.A(cnt_main[4]), .B(cnt_main[2]), .C(cnt_main[3]), 
         .D(cnt_main[0]), .Z(n25800)) /* synthesis lut_function=(A+!(B+(C+(D)))) */ ;
    defparam i1_4_lut_else_4_lut.init = 16'haaab;
    PFUMX mux_131_Mux_0_i18 (.BLUT(n16_adj_5138), .ALUT(n17), .C0(cnt_scan[1]), 
          .Z(n18_adj_5168)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;
    PFUMX i47_adj_251 (.BLUT(n6_adj_5176), .ALUT(n23278), .C0(state[3]), 
          .Z(n24));
    LUT4 i13165_2_lut_rep_461 (.A(cnt_main[3]), .B(cnt_main[2]), .Z(n25743)) /* synthesis lut_function=(A (B)) */ ;
    defparam i13165_2_lut_rep_461.init = 16'h8888;
    LUT4 i1_2_lut_rep_349_3_lut_4_lut (.A(cnt_main[3]), .B(cnt_main[2]), 
         .C(cnt_main[4]), .D(cnt_main[1]), .Z(n25631)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;
    defparam i1_2_lut_rep_349_3_lut_4_lut.init = 16'hf8f0;
    LUT4 i1_2_lut_rep_462 (.A(cnt_main[3]), .B(cnt_main[2]), .Z(n25744)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_462.init = 16'heeee;
    LUT4 equal_8_i9_2_lut_rep_328_3_lut_4_lut (.A(cnt_main[3]), .B(cnt_main[2]), 
         .C(n25750), .D(cnt_main[4]), .Z(n25610)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam equal_8_i9_2_lut_rep_328_3_lut_4_lut.init = 16'hfffe;
    LUT4 i21080_3_lut_3_lut_4_lut_4_lut_4_lut (.A(num2[0]), .B(n25564), 
         .C(n15_adj_5143), .D(n25601), .Z(n23957)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C (D))) */ ;
    defparam i21080_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hf022;
    LUT4 mux_414_Mux_19_i15_3_lut_4_lut_4_lut (.A(num2[0]), .B(n25666), 
         .C(n25635), .D(n25630), .Z(n23761)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B+(C))) */ ;
    defparam mux_414_Mux_19_i15_3_lut_4_lut_4_lut.init = 16'hfc5c;
    LUT4 i21078_3_lut_3_lut_4_lut_4_lut_4_lut (.A(num2[0]), .B(n25564), 
         .C(n15_adj_5120), .D(n25601), .Z(n23955)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C (D))) */ ;
    defparam i21078_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hf022;
    LUT4 i3_4_lut_4_lut (.A(num2[0]), .B(n16320), .C(n5995), .D(cnt_scan[1]), 
         .Z(n20748)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i3_4_lut_4_lut.init = 16'h1000;
    LUT4 n16572_bdd_3_lut_4_lut_4_lut_4_lut (.A(num2[0]), .B(n25564), .C(n16722), 
         .D(n25601), .Z(n25315)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)))+!A (C+!(D)))) */ ;
    defparam n16572_bdd_3_lut_4_lut_4_lut_4_lut.init = 16'h0f22;
    LUT4 n23548_bdd_3_lut (.A(n25586), .B(state[2]), .C(state_back[3]), 
         .Z(n25323)) /* synthesis lut_function=(!(A (B)+!A (B+!(C)))) */ ;
    defparam n23548_bdd_3_lut.init = 16'h3232;
    PFUMX i47_adj_252 (.BLUT(n6_adj_5178), .ALUT(n23279), .C0(state[3]), 
          .Z(n24_adj_5157));
    LUT4 i3_3_lut_4_lut_4_lut_4_lut (.A(num2[0]), .B(n25635), .C(n25601), 
         .D(n25600), .Z(n9_adj_5181)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i3_3_lut_4_lut_4_lut_4_lut.init = 16'h4000;
    LUT4 i5917_4_lut_4_lut (.A(num2[0]), .B(n25753), .C(n25676), .D(cnt_scan[0]), 
         .Z(n8724)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C))+!A (B (C+(D))+!B (C)))) */ ;
    defparam i5917_4_lut_4_lut.init = 16'h21a5;
    LUT4 i17740_2_lut_rep_463 (.A(char[2]), .B(char[1]), .Z(n25745)) /* synthesis lut_function=(A+(B)) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(129[56:62])
    defparam i17740_2_lut_rep_463.init = 16'heeee;
    LUT4 i17745_2_lut_3_lut (.A(char[2]), .B(char[1]), .C(char[3]), .Z(n20442)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(129[56:62])
    defparam i17745_2_lut_3_lut.init = 16'he0e0;
    LUT4 i2_3_lut_rep_389_4_lut (.A(char[2]), .B(char[1]), .C(char[3]), 
         .D(char[4]), .Z(n25671)) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(129[56:62])
    defparam i2_3_lut_rep_389_4_lut.init = 16'he000;
    PFUMX i47_adj_253 (.BLUT(n6_adj_5180), .ALUT(n23281), .C0(state[3]), 
          .Z(n24_adj_5158));
    LUT4 cnt_init_1__bdd_3_lut (.A(cnt_init[1]), .B(cnt_init[2]), .C(n25665), 
         .Z(n26039)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam cnt_init_1__bdd_3_lut.init = 16'h7070;
    LUT4 n1058_bdd_2_lut_22008 (.A(n25324), .B(state[2]), .Z(n25325)) /* synthesis lut_function=(A (B)) */ ;
    defparam n1058_bdd_2_lut_22008.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_adj_254 (.A(cnt_main[0]), .B(cnt_main[1]), .C(cnt_main[4]), 
         .Z(n62_adj_5100)) /* synthesis lut_function=(A (B+(C))+!A ((C)+!B)) */ ;
    defparam i1_2_lut_3_lut_adj_254.init = 16'hf9f9;
    LUT4 i2_2_lut_3_lut (.A(cnt_main[2]), .B(cnt_main[0]), .C(time_data[15]), 
         .Z(n17_adj_5182)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i2_2_lut_3_lut.init = 16'h2020;
    PFUMX i47_adj_255 (.BLUT(n6_adj_5064), .ALUT(n23345), .C0(state[3]), 
          .Z(n26));
    LUT4 i41_1_lut_rep_466 (.A(cnt_scan[4]), .Z(n25748)) /* synthesis lut_function=(!(A)) */ ;
    defparam i41_1_lut_rep_466.init = 16'h5555;
    LUT4 i1_4_lut_4_lut_adj_256 (.A(cnt_scan[4]), .B(n25686), .C(n24908), 
         .D(n25696), .Z(n23310)) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;
    defparam i1_4_lut_4_lut_adj_256.init = 16'hf400;
    PFUMX i22163 (.BLUT(n25784), .ALUT(n25785), .C0(time_data[0]), .Z(n25786));
    LUT4 i20665_2_lut_rep_467 (.A(cnt_main[3]), .B(cnt_main[4]), .Z(n25749)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i20665_2_lut_rep_467.init = 16'hdddd;
    LUT4 i13748_2_lut_3_lut_4_lut (.A(cnt_main[3]), .B(cnt_main[4]), .C(cnt_main[1]), 
         .D(cnt_main[0]), .Z(n15856)) /* synthesis lut_function=((B+(C+!(D)))+!A) */ ;
    defparam i13748_2_lut_3_lut_4_lut.init = 16'hfdff;
    LUT4 i9253_2_lut_3_lut_4_lut_4_lut (.A(n25641), .B(n25605), .C(n2557), 
         .D(n25639), .Z(n12055)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A !(B (D)+!B (C (D))))) */ ;
    defparam i9253_2_lut_3_lut_4_lut_4_lut.init = 16'h7400;
    LUT4 i1_3_lut_4_lut_4_lut (.A(state[3]), .B(state_back[1]), .C(state[0]), 
         .D(state[2]), .Z(n21)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(41[4] 175[11])
    defparam i1_3_lut_4_lut_4_lut.init = 16'h0004;
    LUT4 equal_8_i6_2_lut_rep_468 (.A(cnt_main[0]), .B(cnt_main[1]), .Z(n25750)) /* synthesis lut_function=(A+(B)) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(55[8:12])
    defparam equal_8_i6_2_lut_rep_468.init = 16'heeee;
    PFUMX i30 (.BLUT(n23307), .ALUT(n9_adj_5181), .C0(cnt_scan[1]), .Z(n13_adj_5174));
    LUT4 i13360_2_lut_rep_392_3_lut_4_lut (.A(cnt_main[0]), .B(cnt_main[1]), 
         .C(cnt_main[4]), .D(cnt_main[3]), .Z(n25674)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(55[8:12])
    defparam i13360_2_lut_rep_392_3_lut_4_lut.init = 16'hfeff;
    LUT4 i48_4_lut_4_lut (.A(n25638), .B(state[4]), .C(state_back[4]), 
         .D(state[5]), .Z(n29_adj_5068)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (D)+!B !(C (D))))) */ ;
    defparam i48_4_lut_4_lut.init = 16'h3044;
    PFUMX i21041 (.BLUT(n8_adj_5139), .ALUT(n9_adj_5063), .C0(cnt_scan[1]), 
          .Z(n23918));
    LUT4 i17700_2_lut_rep_470 (.A(char[1]), .B(num2[1]), .Z(n25752)) /* synthesis lut_function=(A+!(B)) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(139[77:83])
    defparam i17700_2_lut_rep_470.init = 16'hbbbb;
    LUT4 i17708_3_lut_4_lut (.A(char[1]), .B(num2[1]), .C(num2[2]), .D(char[2]), 
         .Z(n6_adj_5088)) /* synthesis lut_function=(A ((D)+!C)+!A !(B (C+!(D))+!B !((D)+!C))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(139[77:83])
    defparam i17708_3_lut_4_lut.init = 16'hbf0b;
    LUT4 i13173_3_lut (.A(cnt_main[3]), .B(\tamp_data[7] ), .C(cnt_main[0]), 
         .Z(n80)) /* synthesis lut_function=(!(A+(B (C)))) */ ;
    defparam i13173_3_lut.init = 16'h1515;
    PFUMX i21033 (.BLUT(n11_adj_5131), .ALUT(n12_adj_5053), .C0(cnt_scan[1]), 
          .Z(n23910));
    PFUMX i21039 (.BLUT(n11_adj_5129), .ALUT(n12_adj_5062), .C0(cnt_scan[1]), 
          .Z(n23916));
    PFUMX i22546 (.BLUT(n26493), .ALUT(n23), .C0(state[5]), .Z(n26494));
    LUT4 i2_3_lut_rep_394_4_lut (.A(char[1]), .B(num2[1]), .C(char[2]), 
         .D(num2[2]), .Z(n25676)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(139[77:83])
    defparam i2_3_lut_rep_394_4_lut.init = 16'hb44b;
    PFUMX i21042 (.BLUT(n11_adj_5166), .ALUT(n12_adj_5061), .C0(cnt_scan[1]), 
          .Z(n23919));
    LUT4 i1_4_lut_adj_257 (.A(cnt_main[0]), .B(cnt_main[3]), .C(time_data[17]), 
         .D(time_data[7]), .Z(n102)) /* synthesis lut_function=(!(A ((D)+!B)+!A !(B+!(C)))) */ ;
    defparam i1_4_lut_adj_257.init = 16'h45cd;
    L6MUX21 i21046 (.D0(n23921), .D1(n23922), .SD(cnt_scan[2]), .Z(n23923));
    L6MUX21 i21049 (.D0(n23924), .D1(n23925), .SD(cnt_scan[2]), .Z(n23926));
    PFUMX i4307 (.BLUT(n6104), .ALUT(n7109), .C0(n23861), .Z(n7110));
    LUT4 i1_2_lut_rep_471 (.A(char[1]), .B(num2[1]), .Z(n25753)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut_rep_471.init = 16'h6666;
    LUT4 i3368_3_lut_3_lut_4_lut (.A(char[1]), .B(num2[1]), .C(num2[0]), 
         .D(n25676), .Z(n6170)) /* synthesis lut_function=(!(A (B (D)+!B !(C))+!A !(B (C)+!B !(D)))) */ ;
    defparam i3368_3_lut_3_lut_4_lut.init = 16'h60f9;
    PFUMX i4309 (.BLUT(n8724), .ALUT(n8725), .C0(n25565), .Z(n7112));
    LUT4 i2_4_lut_adj_258 (.A(\tamp_data[9] ), .B(n25764), .C(\tamp_data[5] ), 
         .D(cnt_main[0]), .Z(n32)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i2_4_lut_adj_258.init = 16'hc088;
    LUT4 i1_3_lut_3_lut_4_lut (.A(char[1]), .B(num2[1]), .C(n25676), .D(n25635), 
         .Z(n6178)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam i1_3_lut_3_lut_4_lut.init = 16'h6966;
    LUT4 n9197_bdd_4_lut (.A(n24907), .B(n1355), .C(n31), .D(n1354), 
         .Z(n25411)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A ((D)+!C))) */ ;
    defparam n9197_bdd_4_lut.init = 16'h22f0;
    LUT4 i21523_2_lut_rep_479 (.A(state[2]), .B(state[1]), .Z(n25761)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i21523_2_lut_rep_479.init = 16'h1111;
    PFUMX i21070 (.BLUT(n23945), .ALUT(n23946), .C0(cnt_scan[1]), .Z(n23947));
    PFUMX i22524 (.BLUT(n26454), .ALUT(n26453), .C0(cnt_scan[0]), .Z(n26455));
    LUT4 i2_3_lut_4_lut_adj_259 (.A(char[1]), .B(num2[1]), .C(n25635), 
         .D(n25676), .Z(n6028)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B+(C+(D)))) */ ;
    defparam i2_3_lut_4_lut_adj_259.init = 16'hfff6;
    FD1P3AY oled_rst_369 (.D(n3189[0]), .SP(clk_c_enable_1429), .CK(clk_c), 
            .Q(oled_rst_c)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam oled_rst_369.GSR = "ENABLED";
    PFUMX i22522 (.BLUT(n26450), .ALUT(n26449), .C0(cnt_scan[2]), .Z(n26451));
    LUT4 i3_3_lut_4_lut (.A(n25609), .B(n25692), .C(n20_adj_5102), .D(n42_adj_5155), 
         .Z(clk_c_enable_10)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i3_3_lut_4_lut.init = 16'h1000;
    LUT4 i2_4_lut_4_lut_adj_260 (.A(state[2]), .B(state[0]), .C(state[3]), 
         .D(n25653), .Z(n9_adj_5058)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A (B (C+(D))+!B ((D)+!C)))) */ ;
    defparam i2_4_lut_4_lut_adj_260.init = 16'h0016;
    PFUMX i21079 (.BLUT(n23954), .ALUT(n23955), .C0(cnt_scan[0]), .Z(n23956));
    FD1P3IX cnt_delay_i0_i0 (.D(n2559[0]), .SP(clk_c_enable_1452), .CD(n12055), 
            .CK(clk_c), .Q(cnt_delay[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam cnt_delay_i0_i0.GSR = "ENABLED";
    LUT4 i13903_2_lut_rep_308_3_lut_3_lut_4_lut (.A(char[1]), .B(num2[1]), 
         .C(n25676), .D(num2[0]), .Z(n25590)) /* synthesis lut_function=(!(A (B (C (D)))+!A !(B+!(C (D))))) */ ;
    defparam i13903_2_lut_rep_308_3_lut_3_lut_4_lut.init = 16'h6fff;
    FD1P3IX num2_i0_i0 (.D(num2_7__N_748[0]), .SP(clk_c_enable_1431), .CD(n12049), 
            .CK(clk_c), .Q(num2[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam num2_i0_i0.GSR = "ENABLED";
    FD1P3IX num1_i0_i0 (.D(num1_7__N_732[0]), .SP(clk_c_enable_1432), .CD(n14556), 
            .CK(clk_c), .Q(num1[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam num1_i0_i0.GSR = "ENABLED";
    PFUMX i21082 (.BLUT(n23957), .ALUT(n23958), .C0(cnt_scan[0]), .Z(n23959));
    LUT4 i1_2_lut_3_lut_adj_261 (.A(state[2]), .B(state[1]), .C(state_back[3]), 
         .Z(n8_adj_5183)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_261.init = 16'h1010;
    LUT4 i1_2_lut_rep_282_3_lut_3_lut_4_lut (.A(char[1]), .B(num2[1]), .C(n25676), 
         .D(n25635), .Z(n25564)) /* synthesis lut_function=(A (((D)+!C)+!B)+!A (B+((D)+!C))) */ ;
    defparam i1_2_lut_rep_282_3_lut_3_lut_4_lut.init = 16'hff6f;
    LUT4 i5075_2_lut_rep_293_3_lut_4_lut (.A(char[1]), .B(num2[1]), .C(n25635), 
         .D(n25676), .Z(n25575)) /* synthesis lut_function=(!(A (B+(C (D)+!C !(D)))+!A ((C (D)+!C !(D))+!B))) */ ;
    defparam i5075_2_lut_rep_293_3_lut_4_lut.init = 16'h0660;
    LUT4 i5916_4_lut_4_lut (.A(n25601), .B(n25598), .C(cnt_scan[0]), .D(n6028), 
         .Z(n8723)) /* synthesis lut_function=(A (B+(C))+!A ((D)+!C)) */ ;
    defparam i5916_4_lut_4_lut.init = 16'hfdad;
    LUT4 i1_2_lut_rep_307_3_lut_4_lut (.A(char[1]), .B(num2[1]), .C(n25635), 
         .D(n25676), .Z(n25589)) /* synthesis lut_function=(A ((C+!(D))+!B)+!A (B+(C+!(D)))) */ ;
    defparam i1_2_lut_rep_307_3_lut_4_lut.init = 16'hf6ff;
    LUT4 i20677_2_lut_rep_281_3_lut_3_lut_4_lut (.A(char[1]), .B(num2[1]), 
         .C(n25676), .D(n25635), .Z(n25563)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (((D)+!C)+!B))) */ ;
    defparam i20677_2_lut_rep_281_3_lut_3_lut_4_lut.init = 16'h0060;
    LUT4 equal_1328_i8_2_lut_rep_401_3_lut (.A(state[2]), .B(state[1]), 
         .C(state[0]), .Z(n25683)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam equal_1328_i8_2_lut_rep_401_3_lut.init = 16'hfefe;
    PFUMX i64 (.BLUT(n17_adj_5182), .ALUT(n34_adj_5184), .C0(cnt_main[1]), 
          .Z(n61));
    LUT4 n9339_bdd_4_lut (.A(n25614), .B(state[4]), .C(n25519), .D(cnt_scan[4]), 
         .Z(state_5__N_840[4])) /* synthesis lut_function=(A (C+!(D))+!A (B (C+!(D))+!B (C (D)))) */ ;
    defparam n9339_bdd_4_lut.init = 16'hf0ee;
    LUT4 i9206_3_lut_4_lut_4_lut (.A(n25641), .B(n25604), .C(n25638), 
         .D(n25639), .Z(n12019)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A !(B (D)+!B (C (D))))) */ ;
    defparam i9206_3_lut_4_lut_4_lut.init = 16'h7400;
    LUT4 equal_1334_i8_2_lut_rep_402_3_lut (.A(state[5]), .B(state[4]), 
         .C(state[3]), .Z(n25684)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam equal_1334_i8_2_lut_rep_402_3_lut.init = 16'hfefe;
    LUT4 i2_2_lut_rep_316_3_lut_4_lut (.A(char[1]), .B(num2[1]), .C(n25635), 
         .D(n25676), .Z(n25598)) /* synthesis lut_function=(!(A (B (C (D)))+!A !(B+!(C (D))))) */ ;
    defparam i2_2_lut_rep_316_3_lut_4_lut.init = 16'h6fff;
    LUT4 n25188_bdd_3_lut_4_lut (.A(n23965), .B(cnt_scan[3]), .C(n25187), 
         .D(cnt_scan[4]), .Z(n25189)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C (D))) */ ;
    defparam n25188_bdd_3_lut_4_lut.init = 16'hf088;
    LUT4 n2422_bdd_3_lut_21801_3_lut_4_lut (.A(char[1]), .B(num2[1]), .C(num2[0]), 
         .D(n25676), .Z(n24962)) /* synthesis lut_function=(!(A (B (C)+!B !(D))+!A !(B (D)+!B !(C)))) */ ;
    defparam n2422_bdd_3_lut_21801_3_lut_4_lut.init = 16'h6f09;
    LUT4 n2423_bdd_3_lut_21880_3_lut_4_lut (.A(char[1]), .B(num2[1]), .C(num2[0]), 
         .D(n25676), .Z(n25033)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C (D)+!C !(D)))) */ ;
    defparam n2423_bdd_3_lut_21880_3_lut_4_lut.init = 16'h900f;
    LUT4 i67_4_lut_4_lut (.A(cnt_main[1]), .B(cnt_main[0]), .C(cnt_main[3]), 
         .D(cnt_main[2]), .Z(n65)) /* synthesis lut_function=(A (B (C (D)))+!A !(B+(D))) */ ;
    defparam i67_4_lut_4_lut.init = 16'h8011;
    LUT4 i3193_3_lut_4_lut_4_lut_3_lut_4_lut (.A(char[1]), .B(num2[1]), 
         .C(n25635), .D(n25676), .Z(n5995)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+!(D)))+!A !(B (C+!(D))+!B !((D)+!C)))) */ ;
    defparam i3193_3_lut_4_lut_4_lut_3_lut_4_lut.init = 16'h60f6;
    LUT4 num2_0__bdd_3_lut_3_lut_4_lut (.A(char[1]), .B(num2[1]), .C(num2[0]), 
         .D(n25676), .Z(n23504)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam num2_0__bdd_3_lut_3_lut_4_lut.init = 16'h69f6;
    LUT4 i1_2_lut_3_lut_4_lut_adj_262 (.A(n25760), .B(n25695), .C(n3264), 
         .D(n25691), .Z(n4_adj_5094)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_262.init = 16'he0f0;
    LUT4 i1_2_lut_rep_358_3_lut_4_lut (.A(state[2]), .B(state[1]), .C(state[3]), 
         .D(state[0]), .Z(n25640)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_358_3_lut_4_lut.init = 16'hfffe;
    LUT4 i20684_2_lut_rep_384_3_lut (.A(char[1]), .B(num2[1]), .C(num2[0]), 
         .Z(n25666)) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;
    defparam i20684_2_lut_rep_384_3_lut.init = 16'hf6f6;
    LUT4 i1_4_lut_4_lut_4_lut (.A(n1359), .B(n1358), .C(n25556), .D(num1[0]), 
         .Z(n23378)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A !(B (C)))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(129[51:75])
    defparam i1_4_lut_4_lut_4_lut.init = 16'h6040;
    LUT4 num2_0__bdd_3_lut_21916_3_lut_4_lut (.A(char[1]), .B(num2[1]), 
         .C(num2[0]), .D(n25676), .Z(n14_adj_5119)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)))+!A !(B (C (D))+!B !(C (D)+!C !(D))))) */ ;
    defparam num2_0__bdd_3_lut_21916_3_lut_4_lut.init = 16'h6990;
    LUT4 n2422_bdd_3_lut_22042_4_lut (.A(char[1]), .B(num2[1]), .C(num2[0]), 
         .D(n25676), .Z(n24963)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (D))+!A (B (D)+!B (C (D)+!C !(D))))) */ ;
    defparam n2422_bdd_3_lut_22042_4_lut.init = 16'h09f6;
    PFUMX i21047 (.BLUT(n23360), .ALUT(n9_adj_5052), .C0(cnt_scan[1]), 
          .Z(n23924));
    PFUMX i21038 (.BLUT(n23359), .ALUT(n9_adj_5051), .C0(cnt_scan[1]), 
          .Z(n23915));
    LUT4 i21402_2_lut_rep_480 (.A(cnt_main[1]), .B(cnt_main[0]), .Z(n25762)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i21402_2_lut_rep_480.init = 16'h1111;
    LUT4 equal_1334_i9_2_lut_rep_359_3_lut_3_lut_4_lut (.A(state[5]), .B(state[4]), 
         .C(state[3]), .D(n25761), .Z(n25641)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;
    defparam equal_1334_i9_2_lut_rep_359_3_lut_3_lut_4_lut.init = 16'hfeff;
    PFUMX i32 (.BLUT(n5_adj_5080), .ALUT(n23314), .C0(state[2]), .Z(n15_adj_5071));
    LUT4 i1_2_lut_rep_333_3_lut_4_lut (.A(state[5]), .B(state[4]), .C(state[2]), 
         .D(state[3]), .Z(n25646)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_333_3_lut_4_lut.init = 16'hfffe;
    PFUMX i21045 (.BLUT(n11_adj_5050), .ALUT(n12_adj_5049), .C0(cnt_scan[1]), 
          .Z(n23922));
    LUT4 i13335_4_lut_4_lut (.A(cnt_main[0]), .B(cnt_main[1]), .C(n25718), 
         .D(n25629), .Z(n16111)) /* synthesis lut_function=(A (B+(D))+!A ((C)+!B)) */ ;
    defparam i13335_4_lut_4_lut.init = 16'hfbd9;
    PFUMX i22140 (.BLUT(n25538), .ALUT(n25537), .C0(cnt[3]), .Z(n25539));
    L6MUX21 i21064 (.D0(n23939), .D1(n23940), .SD(cnt_scan[2]), .Z(n23941));
    PFUMX i97 (.BLUT(n69_adj_5173), .ALUT(n23310), .C0(state[3]), .Z(n72));
    LUT4 i21385_2_lut_rep_318_2_lut_4_lut_4_lut (.A(num2[2]), .B(char[2]), 
         .C(char[1]), .D(num2[1]), .Z(n25600)) /* synthesis lut_function=(!(A (B (C+!(D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C+!(D))))) */ ;
    defparam i21385_2_lut_rep_318_2_lut_4_lut_4_lut.init = 16'h0960;
    LUT4 i20927_2_lut_3_lut_3_lut_3_lut_4_lut (.A(char[1]), .B(num2[1]), 
         .C(n25635), .D(n25676), .Z(n23803)) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A ((C+!(D))+!B))) */ ;
    defparam i20927_2_lut_3_lut_3_lut_3_lut_4_lut.init = 16'h0600;
    LUT4 i2_3_lut_4_lut_adj_263 (.A(state[5]), .B(state[4]), .C(state[2]), 
         .D(n17_adj_5171), .Z(n29)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i2_3_lut_4_lut_adj_263.init = 16'h0100;
    LUT4 i1_2_lut_rep_350_4_lut_4_lut (.A(num2[2]), .B(char[2]), .C(char[1]), 
         .D(num2[1]), .Z(n25632)) /* synthesis lut_function=(A (B ((D)+!C)+!B !((D)+!C))+!A !(B ((D)+!C)+!B !((D)+!C))) */ ;
    defparam i1_2_lut_rep_350_4_lut_4_lut.init = 16'h9969;
    PFUMX i21062 (.BLUT(n23379), .ALUT(n9_adj_5047), .C0(cnt_scan[1]), 
          .Z(n23939));
    LUT4 i20842_2_lut_rep_298_3_lut_3_lut_3_lut_4_lut (.A(char[1]), .B(num2[1]), 
         .C(n25635), .D(n25676), .Z(n25580)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C+!(D))+!B (C)))) */ ;
    defparam i20842_2_lut_rep_298_3_lut_3_lut_3_lut_4_lut.init = 16'h0f09;
    PFUMX i21032 (.BLUT(n23378), .ALUT(n9_adj_5046), .C0(cnt_scan[1]), 
          .Z(n23909));
    LUT4 i1_2_lut_4_lut_adj_264 (.A(cnt_init[2]), .B(n25756), .C(cnt_init[0]), 
         .D(state_back[5]), .Z(n19_adj_5179)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (B (D))) */ ;
    defparam i1_2_lut_4_lut_adj_264.init = 16'hec00;
    LUT4 i1_2_lut_3_lut_4_lut_adj_265 (.A(cnt_scan[4]), .B(n25614), .C(n361[6]), 
         .D(state[3]), .Z(n3624[6])) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(111[7] 142[14])
    defparam i1_2_lut_3_lut_4_lut_adj_265.init = 16'h1000;
    LUT4 i43_3_lut_4_lut_3_lut (.A(cnt_main[1]), .B(cnt_main[0]), .C(cnt_main[2]), 
         .Z(n20_adj_5099)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B+!(C)))) */ ;
    defparam i43_3_lut_4_lut_3_lut.init = 16'h1818;
    LUT4 i20848_2_lut_3_lut_4_lut (.A(char[1]), .B(num2[1]), .C(num2[0]), 
         .D(n25676), .Z(n14_adj_5185)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C+!(D)))+!A (B (C+!(D))+!B (C+(D))))) */ ;
    defparam i20848_2_lut_3_lut_4_lut.init = 16'h0609;
    LUT4 i1_2_lut_rep_295_2_lut_3_lut_4_lut (.A(char[1]), .B(num2[1]), .C(n25635), 
         .D(n25676), .Z(n25577)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))) */ ;
    defparam i1_2_lut_rep_295_2_lut_3_lut_4_lut.init = 16'h9669;
    LUT4 i1_2_lut_3_lut_4_lut_adj_266 (.A(cnt_scan[4]), .B(n25614), .C(n361[7]), 
         .D(state[3]), .Z(n3624[7])) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(111[7] 142[14])
    defparam i1_2_lut_3_lut_4_lut_adj_266.init = 16'h1000;
    LUT4 i1_2_lut_rep_348_4_lut_4_lut (.A(num2[2]), .B(char[2]), .C(char[1]), 
         .D(num2[1]), .Z(n25630)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D))))) */ ;
    defparam i1_2_lut_rep_348_4_lut_4_lut.init = 16'h6ff6;
    LUT4 mux_414_Mux_12_i14_4_lut_4_lut_3_lut_4_lut (.A(char[1]), .B(num2[1]), 
         .C(n25676), .D(num2[0]), .Z(n23763)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B !(C+!(D))))) */ ;
    defparam mux_414_Mux_12_i14_4_lut_4_lut_3_lut_4_lut.init = 16'h6f06;
    PFUMX i21048 (.BLUT(n22121), .ALUT(n12_adj_5043), .C0(cnt_scan[1]), 
          .Z(n23925));
    LUT4 i1_4_lut_4_lut_adj_267 (.A(cnt_main[2]), .B(n46), .C(n25762), 
         .D(time_data[1]), .Z(n37)) /* synthesis lut_function=(A (C (D))+!A (B+(C (D)))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(60[8:12])
    defparam i1_4_lut_4_lut_adj_267.init = 16'hf444;
    LUT4 i1_2_lut_4_lut_adj_268 (.A(cnt_init[2]), .B(n25756), .C(cnt_init[0]), 
         .D(state_back[4]), .Z(n19_adj_5177)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (B (D))) */ ;
    defparam i1_2_lut_4_lut_adj_268.init = 16'hec00;
    PFUMX i21063 (.BLUT(n10074), .ALUT(n12_adj_5042), .C0(cnt_scan[1]), 
          .Z(n23940));
    LUT4 i3302_3_lut_3_lut_4_lut (.A(char[1]), .B(num2[1]), .C(n25635), 
         .D(num2[0]), .Z(n6104)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam i3302_3_lut_3_lut_4_lut.init = 16'h6ff0;
    LUT4 i1_2_lut_rep_385_3_lut (.A(char[1]), .B(num2[1]), .C(num2[0]), 
         .Z(n25667)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;
    defparam i1_2_lut_rep_385_3_lut.init = 16'h9696;
    L6MUX21 i21088 (.D0(n23963), .D1(n23964), .SD(cnt_scan[2]), .Z(n23965));
    LUT4 n2423_bdd_2_lut_22046_4_lut_4_lut (.A(num2[2]), .B(char[2]), .C(char[1]), 
         .D(num2[1]), .Z(n25032)) /* synthesis lut_function=(A (B (C+!(D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C+!(D)))) */ ;
    defparam n2423_bdd_2_lut_22046_4_lut_4_lut.init = 16'hf69f;
    LUT4 i1_2_lut_3_lut_4_lut_adj_269 (.A(cnt_scan[4]), .B(n25614), .C(n361[5]), 
         .D(state[3]), .Z(n3624[5])) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(111[7] 142[14])
    defparam i1_2_lut_3_lut_4_lut_adj_269.init = 16'h1000;
    LUT4 i21589_2_lut_2_lut_4_lut_4_lut (.A(num2[2]), .B(char[2]), .C(char[1]), 
         .D(num2[1]), .Z(n23698)) /* synthesis lut_function=(!(A (B+!(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))))) */ ;
    defparam i21589_2_lut_2_lut_4_lut_4_lut.init = 16'h6006;
    LUT4 n15195_bdd_3_lut_22114 (.A(cnt_scan[2]), .B(y_ph[0]), .C(cnt_scan[1]), 
         .Z(n25428)) /* synthesis lut_function=(A (B (C))+!A !(C)) */ ;
    defparam n15195_bdd_3_lut_22114.init = 16'h8585;
    LUT4 i1_3_lut_4_lut_4_lut_4_lut (.A(cnt_main[2]), .B(cnt_main[0]), .C(n25068), 
         .D(cnt_main[4]), .Z(n60)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B (D)+!B ((D)+!C)))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(60[8:12])
    defparam i1_3_lut_4_lut_4_lut_4_lut.init = 16'h00f4;
    LUT4 i2_2_lut_3_lut_4_lut (.A(state[5]), .B(state[4]), .C(n72), .D(state[1]), 
         .Z(clk_c_enable_702)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i2_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i36_3_lut_4_lut_4_lut (.A(cnt_scan[0]), .B(cnt_scan[2]), .C(cnt_scan[1]), 
         .D(cnt_scan[4]), .Z(n16)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A (B+(C+!(D))))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(111[7] 142[14])
    defparam i36_3_lut_4_lut_4_lut.init = 16'h0180;
    LUT4 i1_2_lut_rep_371_3_lut (.A(state[5]), .B(state[4]), .C(state[1]), 
         .Z(n25653)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_371_3_lut.init = 16'hfefe;
    LUT4 n92_bdd_2_lut_4_lut_4_lut (.A(num1[0]), .B(n1359), .C(n1358), 
         .D(n1356), .Z(n24906)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A ((C+(D))+!B))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(129[51:75])
    defparam n92_bdd_2_lut_4_lut_4_lut.init = 16'h0024;
    LUT4 i20732_3_lut_4_lut_4_lut (.A(cnt_main[0]), .B(cnt_main[1]), .C(n25629), 
         .D(cnt_main[2]), .Z(n23589)) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A !(B (C (D))+!B (D)))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(73[29:34])
    defparam i20732_3_lut_4_lut_4_lut.init = 16'h7388;
    LUT4 i1_2_lut_rep_347_3_lut_3_lut (.A(cnt_main[2]), .B(cnt_main[3]), 
         .C(cnt_main[4]), .Z(n25629)) /* synthesis lut_function=(((C)+!B)+!A) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(60[8:12])
    defparam i1_2_lut_rep_347_3_lut_3_lut.init = 16'hf7f7;
    LUT4 mux_414_Mux_13_i7_3_lut_3_lut_3_lut_4_lut_3_lut_4_lut (.A(char[1]), 
         .B(num2[1]), .C(n25676), .D(num2[0]), .Z(n7_adj_5186)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+(D)))+!A (B (C+(D))+!B (C (D)+!C !(D))))) */ ;
    defparam mux_414_Mux_13_i7_3_lut_3_lut_3_lut_4_lut_3_lut_4_lut.init = 16'h0996;
    LUT4 i63_4_lut_then_4_lut (.A(cnt_main[1]), .B(cnt_main[4]), .C(cnt_main[3]), 
         .D(cnt_main[2]), .Z(n25804)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (C+(D)))) */ ;
    defparam i63_4_lut_then_4_lut.init = 16'h2005;
    LUT4 cnt_main_3__bdd_3_lut_22290 (.A(cnt_main[3]), .B(n25871), .C(cnt_main[1]), 
         .Z(n25872)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam cnt_main_3__bdd_3_lut_22290.init = 16'hcaca;
    LUT4 i1_2_lut_rep_376_2_lut (.A(cnt_main[2]), .B(cnt_main[4]), .Z(n25658)) /* synthesis lut_function=((B)+!A) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(60[8:12])
    defparam i1_2_lut_rep_376_2_lut.init = 16'hdddd;
    LUT4 i1_2_lut_4_lut_adj_270 (.A(cnt_init[2]), .B(n25756), .C(cnt_init[0]), 
         .D(state_back[2]), .Z(n19)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (B (D))) */ ;
    defparam i1_2_lut_4_lut_adj_270.init = 16'hec00;
    PFUMX i22111 (.BLUT(n25496), .ALUT(n25495), .C0(state[5]), .Z(n25497));
    LUT4 i1_2_lut_4_lut_adj_271 (.A(cnt_init[2]), .B(n25756), .C(cnt_init[0]), 
         .D(state_back[0]), .Z(n19_adj_5175)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (B (D))) */ ;
    defparam i1_2_lut_4_lut_adj_271.init = 16'hec00;
    LUT4 i1_2_lut_rep_390_2_lut (.A(cnt_main[2]), .B(cnt_main[0]), .Z(n25672)) /* synthesis lut_function=(!(A+!(B))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(60[8:12])
    defparam i1_2_lut_rep_390_2_lut.init = 16'h4444;
    LUT4 i13559_2_lut_rep_472 (.A(state[0]), .B(state[4]), .Z(n25754)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i13559_2_lut_rep_472.init = 16'heeee;
    LUT4 n3_bdd_4_lut_21706_4_lut (.A(cnt_main[2]), .B(\tamp_data[2] ), 
         .C(time_data[6]), .D(cnt_main[1]), .Z(n24713)) /* synthesis lut_function=(!(A+!(B (C+!(D))+!B (C (D))))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(60[8:12])
    defparam n3_bdd_4_lut_21706_4_lut.init = 16'h5044;
    LUT4 cnt_main_3__bdd_4_lut_22291 (.A(cnt_main[3]), .B(cnt_main[2]), 
         .C(cnt_main[4]), .D(cnt_main[0]), .Z(n25871)) /* synthesis lut_function=(!(A (B ((D)+!C))+!A !(B (D)))) */ ;
    defparam cnt_main_3__bdd_4_lut_22291.init = 16'h66a2;
    PFUMX i21086 (.BLUT(n8_adj_5040), .ALUT(n9_adj_5039), .C0(cnt_scan[1]), 
          .Z(n23963));
    LUT4 i20852_2_lut_3_lut_4_lut (.A(state[0]), .B(state[4]), .C(state[2]), 
         .D(state[3]), .Z(n23718)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20852_2_lut_3_lut_4_lut.init = 16'hfffe;
    PFUMX i21044 (.BLUT(n8_adj_5038), .ALUT(n9_adj_5037), .C0(cnt_scan[1]), 
          .Z(n23921));
    LUT4 i1_2_lut_rep_473 (.A(cnt_init[2]), .B(cnt_init[1]), .Z(n25755)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i1_2_lut_rep_473.init = 16'hdddd;
    PFUMX i21087 (.BLUT(n11), .ALUT(n12), .C0(cnt_scan[1]), .Z(n23964));
    LUT4 i1_4_lut_then_4_lut_adj_272 (.A(cnt_main[0]), .B(cnt_main[2]), 
         .C(cnt_main[3]), .D(cnt_main[4]), .Z(n25810)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B ((D)+!C)+!B (C+(D)))) */ ;
    defparam i1_4_lut_then_4_lut_adj_272.init = 16'hffbc;
    LUT4 i1_4_lut_else_4_lut_adj_273 (.A(cnt_main[0]), .B(cnt_main[2]), 
         .C(cnt_main[3]), .D(cnt_main[4]), .Z(n25809)) /* synthesis lut_function=(A (C+(D))+!A ((C+(D))+!B)) */ ;
    defparam i1_4_lut_else_4_lut_adj_273.init = 16'hfff1;
    LUT4 i1_3_lut_3_lut_adj_274 (.A(cnt_main[2]), .B(time_data[19]), .C(cnt_main[0]), 
         .Z(n34_adj_5184)) /* synthesis lut_function=(!(A+!(B+(C)))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(60[8:12])
    defparam i1_3_lut_3_lut_adj_274.init = 16'h5454;
    PFUMX i74 (.BLUT(n34), .ALUT(n41), .C0(state[5]), .Z(n50));
    LUT4 cnt_init_4__I_0_402_i7_2_lut_rep_474 (.A(cnt_init[3]), .B(cnt_init[4]), 
         .Z(n25756)) /* synthesis lut_function=(A+(B)) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(83[8:12])
    defparam cnt_init_4__I_0_402_i7_2_lut_rep_474.init = 16'heeee;
    LUT4 i2_3_lut_rep_368_4_lut (.A(cnt_init[3]), .B(cnt_init[4]), .C(cnt_init[0]), 
         .D(cnt_init[2]), .Z(n25650)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(83[8:12])
    defparam i2_3_lut_rep_368_4_lut.init = 16'hfeee;
    LUT4 i63_4_lut_else_4_lut (.A(cnt_main[1]), .B(cnt_main[4]), .C(cnt_main[3]), 
         .D(cnt_main[2]), .Z(n25803)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i63_4_lut_else_4_lut.init = 16'h2000;
    PFUMX i21002 (.BLUT(n23875), .ALUT(n23876), .C0(cnt_write[2]), .Z(n23879));
    LUT4 i13085_2_lut_rep_481 (.A(cnt_main[2]), .B(cnt_main[4]), .C(cnt_main[3]), 
         .Z(n25763)) /* synthesis lut_function=(A (B+(C))+!A (B+!(C))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(60[8:12])
    defparam i13085_2_lut_rep_481.init = 16'heded;
    LUT4 n12_bdd_4_lut_22117 (.A(n1145), .B(n585), .C(cnt_scan[2]), .D(cnt_scan[3]), 
         .Z(n25430)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !(B (C)+!B (C+(D)))) */ ;
    defparam n12_bdd_4_lut_22117.init = 16'hac0f;
    LUT4 i21486_2_lut_2_lut_4_lut (.A(n25646), .B(state[0]), .C(state[1]), 
         .D(n16632), .Z(n16636)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(51[5:9])
    defparam i21486_2_lut_2_lut_4_lut.init = 16'h0010;
    LUT4 cnt_init_4__I_0_400_i8_2_lut_rep_395_3_lut (.A(cnt_init[3]), .B(cnt_init[4]), 
         .C(cnt_init[2]), .Z(n25677)) /* synthesis lut_function=(A+(B+(C))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(83[8:12])
    defparam cnt_init_4__I_0_400_i8_2_lut_rep_395_3_lut.init = 16'hfefe;
    LUT4 i1_3_lut_4_lut_adj_275 (.A(n25698), .B(n25697), .C(oled_dcn_N_888), 
         .D(state_back[2]), .Z(n9817)) /* synthesis lut_function=(!(A+!(B ((D)+!C)))) */ ;
    defparam i1_3_lut_4_lut_adj_275.init = 16'h4404;
    LUT4 i2_3_lut_4_lut_3_lut_4_lut_4_lut (.A(cnt_main[2]), .B(cnt_main[4]), 
         .C(cnt_main[3]), .D(cnt_main[1]), .Z(n23157)) /* synthesis lut_function=(A (B+(C (D)+!C !(D)))+!A (B+!(C))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(60[8:12])
    defparam i2_3_lut_4_lut_3_lut_4_lut_4_lut.init = 16'hedcf;
    PFUMX mux_414_Mux_13_i15 (.BLUT(n7_adj_5186), .ALUT(n14_adj_5185), .C0(n25635), 
          .Z(n15_adj_5112)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;
    LUT4 i21514_2_lut_rep_346_3_lut_4_lut (.A(cnt_init[3]), .B(cnt_init[4]), 
         .C(cnt_init[0]), .D(cnt_init[2]), .Z(n25628)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(83[8:12])
    defparam i21514_2_lut_rep_346_3_lut_4_lut.init = 16'h0001;
    LUT4 i13197_2_lut_rep_482 (.A(cnt_main[2]), .B(cnt_main[1]), .Z(n25764)) /* synthesis lut_function=(A (B)) */ ;
    defparam i13197_2_lut_rep_482.init = 16'h8888;
    LUT4 i2_2_lut_rep_396_3_lut_4_lut (.A(cnt_init[3]), .B(cnt_init[4]), 
         .C(cnt_init[1]), .D(cnt_init[2]), .Z(n25678)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(83[8:12])
    defparam i2_2_lut_rep_396_3_lut_4_lut.init = 16'hfeff;
    LUT4 i1_2_lut_rep_338_3_lut_4_lut (.A(cnt_init[3]), .B(cnt_init[4]), 
         .C(cnt_init[0]), .D(cnt_init[2]), .Z(n25620)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(83[8:12])
    defparam i1_2_lut_rep_338_3_lut_4_lut.init = 16'h0010;
    LUT4 cnt_scan_0__bdd_4_lut_22034 (.A(cnt_scan[0]), .B(n23504), .C(num2[0]), 
         .D(n25630), .Z(n25372)) /* synthesis lut_function=(!(A (C+(D))+!A !(B))) */ ;
    defparam cnt_scan_0__bdd_4_lut_22034.init = 16'h444e;
    LUT4 cnt_scan_0__bdd_4_lut_22638 (.A(cnt_scan[0]), .B(n25676), .C(num2[0]), 
         .D(n25753), .Z(n25373)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A !(B ((D)+!C)+!B !(C))) */ ;
    defparam cnt_scan_0__bdd_4_lut_22638.init = 16'h9872;
    LUT4 i1_2_lut_rep_277_3_lut_4_lut (.A(n25698), .B(n25697), .C(n25755), 
         .D(oled_dcn_N_888), .Z(n25559)) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B (C))) */ ;
    defparam i1_2_lut_rep_277_3_lut_4_lut.init = 16'hf4f0;
    PFUMX i22098 (.BLUT(n25470), .ALUT(n25469), .C0(n3599), .Z(cnt_scan_4__N_682[4]));
    LUT4 i1_3_lut_4_lut_adj_276 (.A(cnt_scan[0]), .B(n25566), .C(n1358), 
         .D(num1[0]), .Z(n23379)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))) */ ;
    defparam i1_3_lut_4_lut_adj_276.init = 16'h8008;
    PFUMX i10774 (.BLUT(n13577), .ALUT(n21246), .C0(oled_dcn_N_888), .Z(n13581));
    LUT4 i2718_2_lut_rep_476 (.A(cnt_write[1]), .B(cnt_write[0]), .Z(n25758)) /* synthesis lut_function=(A (B)) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(146[25:41])
    defparam i2718_2_lut_rep_476.init = 16'h8888;
    LUT4 i1_2_lut_4_lut_adj_277 (.A(cnt_scan[0]), .B(n25622), .C(n25566), 
         .D(num1[0]), .Z(n23359)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_4_lut_adj_277.init = 16'h8000;
    LUT4 i1_3_lut_rep_375_4_lut (.A(cnt_main[2]), .B(cnt_main[1]), .C(cnt_main[3]), 
         .D(cnt_main[4]), .Z(n25657)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A ((D)+!C))) */ ;
    defparam i1_3_lut_rep_375_4_lut.init = 16'h0078;
    CCU2D sub_79_add_2_9 (.A0(num1[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n20526), 
          .S0(n361[7]));   // g:/fpga/mxo2/system/project/oled12832.v(121[49:60])
    defparam sub_79_add_2_9.INIT0 = 16'h5555;
    defparam sub_79_add_2_9.INIT1 = 16'h0000;
    defparam sub_79_add_2_9.INJECT1_0 = "NO";
    defparam sub_79_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_79_add_2_7 (.A0(num1[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(num1[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n20525), 
          .COUT(n20526), .S0(n361[5]), .S1(n361[6]));   // g:/fpga/mxo2/system/project/oled12832.v(121[49:60])
    defparam sub_79_add_2_7.INIT0 = 16'h5555;
    defparam sub_79_add_2_7.INIT1 = 16'h5555;
    defparam sub_79_add_2_7.INJECT1_0 = "NO";
    defparam sub_79_add_2_7.INJECT1_1 = "NO";
    LUT4 i2723_2_lut_3_lut (.A(cnt_write[1]), .B(cnt_write[0]), .C(cnt_write[2]), 
         .Z(n2535[2])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(146[25:41])
    defparam i2723_2_lut_3_lut.init = 16'h7878;
    FD1P3IX cnt_write_i0_i0 (.D(n4_adj_5126), .SP(clk_c_enable_1436), .CD(n12019), 
            .CK(clk_c), .Q(cnt_write[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam cnt_write_i0_i0.GSR = "ENABLED";
    PFUMX i21003 (.BLUT(n23877), .ALUT(n23878), .C0(cnt_write[2]), .Z(n23880));
    PFUMX i46 (.BLUT(n5), .ALUT(n8_adj_5183), .C0(state[5]), .Z(n23_adj_5070));
    LUT4 i6068_3_lut (.A(cnt_scan[3]), .B(n322), .C(cnt_scan[0]), .Z(n8876)) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)))) */ ;
    defparam i6068_3_lut.init = 16'h3535;
    CCU2D sub_79_add_2_5 (.A0(num1[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(num1[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n20524), 
          .COUT(n20525), .S0(num1_7__N_732[3]), .S1(num1_7__N_732[4]));   // g:/fpga/mxo2/system/project/oled12832.v(121[49:60])
    defparam sub_79_add_2_5.INIT0 = 16'h5555;
    defparam sub_79_add_2_5.INIT1 = 16'h5555;
    defparam sub_79_add_2_5.INJECT1_0 = "NO";
    defparam sub_79_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_79_add_2_3 (.A0(num1[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(num1[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n20523), 
          .COUT(n20524), .S0(num1_7__N_732[1]), .S1(num1_7__N_732[2]));   // g:/fpga/mxo2/system/project/oled12832.v(121[49:60])
    defparam sub_79_add_2_3.INIT0 = 16'h5555;
    defparam sub_79_add_2_3.INIT1 = 16'h5555;
    defparam sub_79_add_2_3.INJECT1_0 = "NO";
    defparam sub_79_add_2_3.INJECT1_1 = "NO";
    LUT4 i2_3_lut_4_lut_adj_278 (.A(state[1]), .B(n25760), .C(n23590), 
         .D(state[3]), .Z(n27_adj_5133)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i2_3_lut_4_lut_adj_278.init = 16'hfffe;
    CCU2D sub_79_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(num1[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n20523), 
          .S1(num1_7__N_732[0]));   // g:/fpga/mxo2/system/project/oled12832.v(121[49:60])
    defparam sub_79_add_2_1.INIT0 = 16'hF000;
    defparam sub_79_add_2_1.INIT1 = 16'h5555;
    defparam sub_79_add_2_1.INJECT1_0 = "NO";
    defparam sub_79_add_2_1.INJECT1_1 = "NO";
    PFUMX i22188 (.BLUT(n25821), .ALUT(n25822), .C0(state[1]), .Z(n25823));
    LUT4 i21001_3_lut (.A(char_reg[4]), .B(char_reg[0]), .C(cnt_write[3]), 
         .Z(n23878)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21001_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_279 (.A(state[5]), .B(state[4]), .C(state[1]), 
         .D(state[3]), .Z(n16443)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_279.init = 16'hfffe;
    LUT4 state_1__bdd_4_lut_then_4_lut (.A(cnt_scan[0]), .B(cnt_scan[1]), 
         .C(cnt_scan[2]), .D(cnt_scan[3]), .Z(n25822)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A ((C+!(D))+!B))) */ ;
    defparam state_1__bdd_4_lut_then_4_lut.init = 16'h0402;
    FD1P3IX cnt_delay_i0_i15 (.D(n2559[15]), .SP(clk_c_enable_1452), .CD(n12055), 
            .CK(clk_c), .Q(cnt_delay[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam cnt_delay_i0_i15.GSR = "ENABLED";
    FD1P3IX cnt_delay_i0_i14 (.D(n2559[14]), .SP(clk_c_enable_1452), .CD(n12055), 
            .CK(clk_c), .Q(cnt_delay[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam cnt_delay_i0_i14.GSR = "ENABLED";
    FD1P3IX cnt_delay_i0_i13 (.D(n2559[13]), .SP(clk_c_enable_1452), .CD(n12055), 
            .CK(clk_c), .Q(cnt_delay[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam cnt_delay_i0_i13.GSR = "ENABLED";
    FD1P3IX cnt_delay_i0_i12 (.D(n2559[12]), .SP(clk_c_enable_1452), .CD(n12055), 
            .CK(clk_c), .Q(cnt_delay[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam cnt_delay_i0_i12.GSR = "ENABLED";
    FD1P3IX cnt_delay_i0_i11 (.D(n2559[11]), .SP(clk_c_enable_1452), .CD(n12055), 
            .CK(clk_c), .Q(cnt_delay[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam cnt_delay_i0_i11.GSR = "ENABLED";
    PFUMX mux_1283_i4 (.BLUT(n331[3]), .ALUT(n8876), .C0(n3599), .Z(cnt_scan_4__N_682[3]));
    LUT4 n15195_bdd_2_lut_22113_4_lut (.A(n725), .B(n1285), .C(cnt_scan[2]), 
         .D(cnt_scan[1]), .Z(n25427)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(27[33:41])
    defparam n15195_bdd_2_lut_22113_4_lut.init = 16'hca00;
    LUT4 state_1__bdd_4_lut_else_4_lut (.A(cnt_scan[0]), .B(cnt_scan[1]), 
         .C(cnt_scan[2]), .D(cnt_scan[3]), .Z(n25821)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam state_1__bdd_4_lut_else_4_lut.init = 16'h0400;
    L6MUX21 i22073 (.D0(n25431), .D1(n25429), .SD(cnt_scan[0]), .Z(n23935));
    CCU2D sub_104_add_2_9 (.A0(num2[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n20522), 
          .S0(num2_7__N_748[7]));   // g:/fpga/mxo2/system/project/oled12832.v(131[50:61])
    defparam sub_104_add_2_9.INIT0 = 16'h5555;
    defparam sub_104_add_2_9.INIT1 = 16'h0000;
    defparam sub_104_add_2_9.INJECT1_0 = "NO";
    defparam sub_104_add_2_9.INJECT1_1 = "NO";
    PFUMX i22071 (.BLUT(n12_adj_5045), .ALUT(n25430), .C0(cnt_scan[1]), 
          .Z(n25431));
    LUT4 i2730_2_lut_3_lut_4_lut (.A(cnt_write[1]), .B(cnt_write[0]), .C(cnt_write[3]), 
         .D(cnt_write[2]), .Z(n2535[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(146[25:41])
    defparam i2730_2_lut_3_lut_4_lut.init = 16'h78f0;
    CCU2D sub_104_add_2_7 (.A0(num2[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(num2[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n20521), 
          .COUT(n20522), .S0(num2_7__N_748[5]), .S1(num2_7__N_748[6]));   // g:/fpga/mxo2/system/project/oled12832.v(131[50:61])
    defparam sub_104_add_2_7.INIT0 = 16'h5555;
    defparam sub_104_add_2_7.INIT1 = 16'h5555;
    defparam sub_104_add_2_7.INJECT1_0 = "NO";
    defparam sub_104_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_104_add_2_5 (.A0(num2[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(num2[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n20520), 
          .COUT(n20521), .S0(num2_7__N_748[3]), .S1(num2_7__N_748[4]));   // g:/fpga/mxo2/system/project/oled12832.v(131[50:61])
    defparam sub_104_add_2_5.INIT0 = 16'h5555;
    defparam sub_104_add_2_5.INIT1 = 16'h5555;
    defparam sub_104_add_2_5.INJECT1_0 = "NO";
    defparam sub_104_add_2_5.INJECT1_1 = "NO";
    FD1P3IX cnt_delay_i0_i10 (.D(n2559[10]), .SP(clk_c_enable_1452), .CD(n12055), 
            .CK(clk_c), .Q(cnt_delay[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam cnt_delay_i0_i10.GSR = "ENABLED";
    PFUMX i22180 (.BLUT(n25809), .ALUT(n25810), .C0(cnt_main[1]), .Z(n16743));
    FD1P3AX cnt_scan_i0_i2 (.D(n21243), .SP(clk_c_enable_1446), .CK(clk_c), 
            .Q(cnt_scan[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam cnt_scan_i0_i2.GSR = "ENABLED";
    PFUMX i22069 (.BLUT(n25428), .ALUT(n25427), .C0(cnt_scan[3]), .Z(n25429));
    PFUMX i22176 (.BLUT(n25803), .ALUT(n25804), .C0(char[6]), .Z(n25805));
    FD1P3IX cnt_delay_i0_i9 (.D(n2559[9]), .SP(clk_c_enable_1452), .CD(n12055), 
            .CK(clk_c), .Q(cnt_delay[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam cnt_delay_i0_i9.GSR = "ENABLED";
    FD1P3IX cnt_delay_i0_i8 (.D(n2559[8]), .SP(clk_c_enable_1452), .CD(n12055), 
            .CK(clk_c), .Q(cnt_delay[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam cnt_delay_i0_i8.GSR = "ENABLED";
    FD1P3IX cnt_delay_i0_i7 (.D(n2559[7]), .SP(clk_c_enable_1452), .CD(n12055), 
            .CK(clk_c), .Q(cnt_delay[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam cnt_delay_i0_i7.GSR = "ENABLED";
    CCU2D sub_104_add_2_3 (.A0(num2[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(num2[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n20519), 
          .COUT(n20520), .S0(num2_7__N_748[1]), .S1(num2_7__N_748[2]));   // g:/fpga/mxo2/system/project/oled12832.v(131[50:61])
    defparam sub_104_add_2_3.INIT0 = 16'h5555;
    defparam sub_104_add_2_3.INIT1 = 16'h5555;
    defparam sub_104_add_2_3.INJECT1_0 = "NO";
    defparam sub_104_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_104_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(num2[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n20519), 
          .S1(num2_7__N_748[0]));   // g:/fpga/mxo2/system/project/oled12832.v(131[50:61])
    defparam sub_104_add_2_1.INIT0 = 16'hF000;
    defparam sub_104_add_2_1.INIT1 = 16'h5555;
    defparam sub_104_add_2_1.INJECT1_0 = "NO";
    defparam sub_104_add_2_1.INJECT1_1 = "NO";
    FD1P3IX cnt_delay_i0_i6 (.D(n2559[6]), .SP(clk_c_enable_1452), .CD(n12055), 
            .CK(clk_c), .Q(cnt_delay[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam cnt_delay_i0_i6.GSR = "ENABLED";
    LUT4 mux_3021_i2_4_lut (.A(n9), .B(n5817[0]), .C(n25587), .D(n16666), 
         .Z(n5820[1])) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam mux_3021_i2_4_lut.init = 16'hc5c0;
    LUT4 n9197_bdd_4_lut_22058 (.A(n25566), .B(n1358), .C(n1359), .D(num1[0]), 
         .Z(n25410)) /* synthesis lut_function=(!((B (C)+!B (C+!(D)))+!A)) */ ;
    defparam n9197_bdd_4_lut_22058.init = 16'h0a08;
    LUT4 i1849_2_lut_rep_477 (.A(cnt_init[0]), .B(cnt_init[1]), .Z(n25759)) /* synthesis lut_function=(A (B)) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(41[4] 175[11])
    defparam i1849_2_lut_rep_477.init = 16'h8888;
    LUT4 i2658_2_lut_3_lut_4_lut (.A(cnt_init[0]), .B(cnt_init[1]), .C(cnt_init[3]), 
         .D(cnt_init[2]), .Z(n1[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // g:/fpga/mxo2/system/project/oled12832.v(41[4] 175[11])
    defparam i2658_2_lut_3_lut_4_lut.init = 16'h78f0;
    PFUMX i22059 (.BLUT(n25411), .ALUT(n25410), .C0(cnt_scan[0]), .Z(n25412));
    FD1P3IX cnt_delay_i0_i5 (.D(n2559[5]), .SP(clk_c_enable_1452), .CD(n12055), 
            .CK(clk_c), .Q(cnt_delay[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=11, LSE_RCOL=2, LSE_LLINE=70, LSE_RLINE=80 */ ;   // g:/fpga/mxo2/system/project/oled12832.v(40[12] 176[6])
    defparam cnt_delay_i0_i5.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module beeper_control
//

module beeper_control (\data_buffer[538] , n26793, \data_buffer[539] , 
            \data_buffer[540] , \data_buffer[544] , \data_buffer[545] , 
            \data_buffer[546] , \data_buffer[547] , \data_buffer[548] , 
            \data_buffer[552] , \data_buffer[553] , \data_buffer[554] , 
            \data_buffer[555] , \data_buffer[556] , \data_buffer[560] , 
            \data_buffer[561] , \data_buffer[562] , \data_buffer[563] , 
            \data_buffer[564] , \data_buffer[568] , \data_buffer[160] , 
            \data_buffer[569] , \data_buffer[570] , \data_buffer[571] , 
            clk_c, \data_buffer[572] , \data_buffer[576] , \data_buffer[577] , 
            \data_buffer[416] , \data_buffer[578] , \data_buffer[579] , 
            \data_buffer[580] , \data_buffer[584] , \data_buffer[585] , 
            \data_buffer[586] , \data_buffer[587] , \data_buffer[588] , 
            \data_buffer[592] , \data_buffer[593] , \data_buffer[594] , 
            \data_buffer[595] , \data_buffer[596] , \data_buffer[600] , 
            \data_buffer[601] , \data_buffer[602] , \data_buffer[603] , 
            \data_buffer[604] , \data_buffer[608] , \data_buffer[609] , 
            \data_buffer[610] , \data_buffer[611] , \data_buffer[612] , 
            \data_buffer[616] , \data_buffer[617] , \data_buffer[618] , 
            \data_buffer[619] , \data_buffer[620] , \data_buffer[624] , 
            \data_buffer[625] , \data_buffer[626] , \data_buffer[627] , 
            \data_buffer[628] , data_length_reg, n15, \data_buffer[632] , 
            \data_buffer[633] , \data_buffer[634] , \data_buffer[635] , 
            \data_buffer[636] , \data_buffer[640] , \data_buffer[641] , 
            \data_buffer[642] , \data_buffer[643] , \data_buffer[644] , 
            \data_buffer[648] , \data_buffer[649] , \data_buffer[650] , 
            \data_buffer[651] , \data_buffer[652] , \data_buffer[656] , 
            \data_buffer[657] , \data_buffer[658] , \data_buffer[659] , 
            \data_buffer[660] , \data_buffer[664] , \data_buffer[665] , 
            \data_buffer[666] , \data_buffer[667] , \data_buffer[668] , 
            \data_buffer[672] , \data_buffer[673] , \data_buffer[674] , 
            \data_buffer[675] , \data_buffer[676] , \data_buffer[680] , 
            \data_buffer[681] , \data_buffer[682] , \data_buffer[683] , 
            \data_buffer[684] , \data_buffer[688] , \data_buffer[689] , 
            \data_buffer[690] , \data_buffer[691] , \data_buffer[692] , 
            \data_buffer[696] , \data_buffer[697] , \data_buffer[698] , 
            \data_buffer[699] , \data_buffer[700] , \data_buffer[704] , 
            \data_buffer[705] , \data_buffer[706] , \data_buffer[707] , 
            \data_buffer[708] , \data_buffer[712] , \data_buffer[713] , 
            \data_buffer[714] , \data_buffer[715] , \data_buffer[716] , 
            \data_buffer[720] , \data_buffer[161] , \data_buffer[721] , 
            \data_buffer[722] , \data_buffer[723] , \data_buffer[724] , 
            \data_buffer[728] , \data_buffer[729] , \data_buffer[730] , 
            \data_buffer[731] , \data_buffer[732] , \data_buffer[736] , 
            \data_buffer[737] , \data_buffer[162] , \data_buffer[738] , 
            \data_buffer[739] , \data_buffer[740] , \data_buffer[744] , 
            \data_buffer[163] , \data_buffer[745] , \data_buffer[746] , 
            \data_buffer[747] , \data_buffer[748] , \data_buffer[752] , 
            \data_buffer[753] , \data_buffer[754] , \data_buffer[755] , 
            \data_buffer[756] , \data_buffer[760] , \data_buffer[761] , 
            \data_buffer[762] , \data_buffer[763] , \data_buffer[764] , 
            \data_buffer[768] , \data_buffer[769] , \data_buffer[770] , 
            \data_buffer[771] , \data_buffer[772] , \data_buffer[776] , 
            \data_buffer[777] , \data_buffer[778] , \data_buffer[779] , 
            \data_buffer[780] , \data_buffer[784] , \data_buffer[785] , 
            \data_buffer[786] , \data_buffer[787] , \data_buffer[788] , 
            \data_buffer[792] , \data_buffer[793] , \data_buffer[794] , 
            \data_buffer[164] , \data_buffer[795] , \data_buffer[796] , 
            \data_buffer[800] , \data_buffer[801] , \data_buffer[802] , 
            \data_buffer[803] , \data_buffer[804] , \data_buffer[808] , 
            \data_buffer[809] , \data_buffer[810] , \data_buffer[811] , 
            \data_buffer[812] , \data_buffer[816] , \data_buffer[817] , 
            \data_buffer[818] , \data_buffer[819] , \data_buffer[820] , 
            \data_buffer[824] , \data_buffer[825] , \data_buffer[826] , 
            \data_buffer[827] , \data_buffer[828] , \data_buffer[832] , 
            \data_buffer[833] , \data_buffer[834] , \data_buffer[835] , 
            \data_buffer[836] , \data_buffer[840] , \data_buffer[841] , 
            \data_buffer[842] , \data_buffer[843] , \data_buffer[844] , 
            \data_buffer[848] , \data_buffer[849] , \data_buffer[850] , 
            \data_buffer[851] , \data_buffer[852] , \data_buffer[856] , 
            \data_buffer[857] , \data_buffer[858] , \data_buffer[859] , 
            \data_buffer[860] , \data_buffer[864] , \data_buffer[865] , 
            \data_buffer[866] , \data_buffer[867] , \data_buffer[868] , 
            \data_buffer[872] , \data_buffer[873] , \data_buffer[874] , 
            \data_buffer[875] , \data_buffer[876] , \data_buffer[880] , 
            \data_buffer[881] , \data_buffer[882] , \data_buffer[883] , 
            \data_buffer[884] , \data_buffer[888] , \data_buffer[889] , 
            \data_buffer[890] , \data_buffer[891] , \data_buffer[892] , 
            \data_buffer[386] , \data_buffer[896] , \data_buffer[897] , 
            \data_buffer[898] , \data_buffer[899] , \data_buffer[900] , 
            \data_buffer[904] , \data_buffer[905] , \data_buffer[906] , 
            \data_buffer[907] , \data_buffer[908] , \data_buffer[912] , 
            \data_buffer[913] , \data_buffer[914] , \data_buffer[915] , 
            \data_buffer[916] , \data_buffer[920] , \data_buffer[921] , 
            \data_buffer[922] , \data_buffer[923] , \data_buffer[924] , 
            \data_buffer[928] , \data_buffer[929] , \data_buffer[930] , 
            \data_buffer[931] , \data_buffer[932] , \data_buffer[168] , 
            \data_buffer[936] , \data_buffer[937] , \data_buffer[938] , 
            \data_buffer[939] , \data_buffer[940] , \data_buffer[944] , 
            \data_buffer[945] , \data_buffer[946] , \data_buffer[947] , 
            \data_buffer[948] , \data_buffer[169] , \data_buffer[170] , 
            \data_buffer[171] , \data_buffer[0] , \data_buffer[387] , 
            \data_buffer[172] , \data_buffer[176] , \data_buffer[177] , 
            \data_buffer[178] , \data_buffer[956] , \data_buffer[179] , 
            \data_buffer[1] , \data_buffer[2] , \data_buffer[3] , \data_buffer[4] , 
            \data_buffer[8] , \data_buffer[9] , \data_buffer[10] , \data_buffer[11] , 
            \data_buffer[12] , \data_buffer[16] , \data_buffer[17] , \data_buffer[18] , 
            \data_buffer[19] , \data_buffer[20] , \data_buffer[24] , \data_buffer[25] , 
            \data_buffer[26] , \data_buffer[27] , \data_buffer[28] , \data_buffer[32] , 
            \data_buffer[33] , \data_buffer[955] , \data_buffer[34] , 
            \data_buffer[35] , \data_buffer[36] , \data_buffer[40] , \data_buffer[41] , 
            \data_buffer[42] , \data_buffer[43] , \data_buffer[44] , \data_buffer[48] , 
            \data_buffer[49] , \data_buffer[50] , \data_buffer[51] , \data_buffer[52] , 
            \data_buffer[56] , \data_buffer[57] , \data_buffer[58] , \data_buffer[954] , 
            \data_buffer[59] , \data_buffer[60] , \data_buffer[388] , 
            \data_buffer[64] , \data_buffer[953] , \data_buffer[952] , 
            \data_buffer[65] , \data_buffer[180] , \data_buffer[66] , 
            \data_buffer[67] , \data_buffer[68] , \data_buffer[72] , \data_buffer[73] , 
            \data_buffer[74] , \data_buffer[75] , \data_buffer[76] , \data_buffer[80] , 
            \data_buffer[81] , \data_buffer[82] , \data_buffer[83] , \data_buffer[84] , 
            \data_buffer[88] , \data_buffer[184] , \data_buffer[89] , 
            \data_buffer[90] , \data_buffer[185] , \data_buffer[91] , 
            \data_buffer[92] , \data_buffer[96] , \data_buffer[97] , \data_buffer[98] , 
            \data_buffer[99] , \data_buffer[100] , \data_buffer[186] , 
            \data_buffer[104] , \data_buffer[105] , \data_buffer[106] , 
            \data_buffer[107] , \data_buffer[108] , \data_buffer[112] , 
            \data_buffer[113] , \data_buffer[114] , \data_buffer[115] , 
            \data_buffer[116] , \data_buffer[120] , \data_buffer[121] , 
            \data_buffer[122] , \data_buffer[123] , \data_buffer[124] , 
            \data_buffer[128] , \data_buffer[129] , \data_buffer[187] , 
            \data_buffer[130] , \data_buffer[131] , \data_buffer[132] , 
            \data_buffer[136] , \data_buffer[137] , \data_buffer[138] , 
            \data_buffer[139] , \data_buffer[140] , \data_buffer[144] , 
            \data_buffer[145] , \data_buffer[146] , \data_buffer[147] , 
            \data_buffer[148] , \data_buffer[152] , \data_buffer[153] , 
            \data_buffer[154] , \data_buffer[155] , \data_buffer[156] , 
            \data_buffer[188] , \data_buffer[392] , \data_buffer[393] , 
            \data_buffer[394] , \data_buffer[192] , \data_buffer[193] , 
            \data_buffer[194] , \data_buffer[195] , \data_buffer[196] , 
            \data_buffer[200] , \data_buffer[395] , \data_buffer[396] , 
            \data_buffer[201] , \data_buffer[202] , \data_buffer[203] , 
            \data_buffer[204] , \data_buffer[208] , \data_buffer[417] , 
            \data_buffer[418] , \data_buffer[419] , \data_buffer[420] , 
            \data_buffer[400] , \data_buffer[401] , \data_buffer[209] , 
            \data_buffer[210] , \data_buffer[424] , \data_buffer[211] , 
            \data_buffer[425] , \data_buffer[212] , \data_buffer[426] , 
            \data_buffer[402] , \data_buffer[427] , \data_buffer[428] , 
            \data_buffer[216] , \data_buffer[217] , \data_buffer[218] , 
            \data_buffer[219] , \data_buffer[432] , \data_buffer[433] , 
            \data_buffer[220] , \data_buffer[434] , \data_buffer[435] , 
            \data_buffer[436] , \data_buffer[440] , \data_buffer[224] , 
            \data_buffer[225] , \data_buffer[441] , \data_buffer[403] , 
            \data_buffer[226] , \data_buffer[227] , \data_buffer[228] , 
            \data_buffer[232] , \data_buffer[233] , \data_buffer[234] , 
            \data_buffer[442] , \data_buffer[443] , \data_buffer[404] , 
            \data_buffer[444] , \data_buffer[235] , \data_buffer[236] , 
            \data_buffer[408] , \data_buffer[240] , \data_buffer[409] , 
            \data_buffer[241] , \data_buffer[448] , \data_buffer[242] , 
            \data_buffer[449] , \data_buffer[450] , \data_buffer[243] , 
            \data_buffer[451] , \data_buffer[244] , \data_buffer[248] , 
            \data_buffer[452] , \data_buffer[249] , \data_buffer[250] , 
            \data_buffer[251] , \data_buffer[252] , \data_buffer[256] , 
            \data_buffer[257] , \data_buffer[258] , \data_buffer[259] , 
            \data_buffer[260] , \data_buffer[264] , \data_buffer[265] , 
            \data_buffer[266] , \data_buffer[267] , \data_buffer[268] , 
            \data_buffer[272] , \data_buffer[456] , \data_buffer[273] , 
            \data_buffer[274] , \data_buffer[457] , \data_buffer[275] , 
            \data_buffer[276] , \data_buffer[458] , data_length, GND_net, 
            \data_buffer[280] , \data_buffer[459] , \data_buffer[460] , 
            \data_buffer[281] , \data_buffer[282] , \data_buffer[283] , 
            \data_buffer[284] , \data_buffer[288] , \data_buffer[464] , 
            \data_buffer[289] , \data_buffer[465] , \data_buffer[290] , 
            \data_buffer[466] , \data_buffer[291] , \data_buffer[292] , 
            \data_buffer[296] , \data_buffer[467] , \data_buffer[297] , 
            \data_buffer[298] , \data_buffer[468] , \data_buffer[472] , 
            \data_buffer[299] , \data_buffer[300] , \data_buffer[304] , 
            \data_buffer[305] , \data_buffer[306] , \data_buffer[307] , 
            \data_buffer[308] , \data_buffer[312] , \data_buffer[473] , 
            \data_buffer[313] , \data_buffer[314] , \data_buffer[315] , 
            \data_buffer[474] , \data_buffer[316] , \data_buffer[475] , 
            \data_buffer[320] , \data_buffer[321] , \data_buffer[476] , 
            \data_buffer[480] , \data_buffer[322] , \data_buffer[323] , 
            \data_buffer[324] , \data_buffer[481] , \data_buffer[328] , 
            \data_buffer[329] , \data_buffer[330] , \data_buffer[331] , 
            \data_buffer[482] , \data_buffer[483] , \data_buffer[484] , 
            \data_buffer[332] , \data_buffer[488] , \data_buffer[336] , 
            \data_buffer[337] , \data_buffer[489] , \data_buffer[338] , 
            \data_buffer[490] , \data_buffer[339] , \data_buffer[491] , 
            \data_buffer[340] , \data_buffer[344] , \data_buffer[492] , 
            \data_buffer[345] , \data_buffer[496] , \data_buffer[497] , 
            \data_buffer[346] , \data_buffer[347] , \data_buffer[498] , 
            \data_buffer[499] , \data_buffer[500] , \data_buffer[348] , 
            \data_buffer[352] , \data_buffer[353] , \data_buffer[354] , 
            \data_buffer[355] , \data_buffer[356] , \data_buffer[504] , 
            \data_buffer[360] , \data_buffer[361] , \data_buffer[505] , 
            \data_buffer[506] , \data_buffer[362] , \data_buffer[507] , 
            \data_buffer[363] , \data_buffer[508] , \data_buffer[364] , 
            \data_buffer[368] , \data_buffer[369] , \data_buffer[512] , 
            \data_buffer[513] , \data_buffer[514] , \data_buffer[515] , 
            \data_buffer[370] , \data_buffer[516] , \data_buffer[520] , 
            \data_buffer[371] , \data_buffer[521] , \data_buffer[372] , 
            \data_buffer[522] , \data_buffer[523] , \data_buffer[524] , 
            \data_buffer[376] , \data_buffer[528] , \data_buffer[529] , 
            \data_buffer[530] , \data_buffer[531] , \data_buffer[532] , 
            \data_buffer[536] , \data_buffer[537] , \data_buffer[377] , 
            \data_buffer[378] , \data_buffer[379] , \data_buffer[380] , 
            \data_buffer[410] , \data_buffer[411] , \data_buffer[412] , 
            \data_buffer[384] , \data_buffer[385] , piano_out_c) /* synthesis syn_module_defined=1 */ ;
    input \data_buffer[538] ;
    input n26793;
    input \data_buffer[539] ;
    input \data_buffer[540] ;
    input \data_buffer[544] ;
    input \data_buffer[545] ;
    input \data_buffer[546] ;
    input \data_buffer[547] ;
    input \data_buffer[548] ;
    input \data_buffer[552] ;
    input \data_buffer[553] ;
    input \data_buffer[554] ;
    input \data_buffer[555] ;
    input \data_buffer[556] ;
    input \data_buffer[560] ;
    input \data_buffer[561] ;
    input \data_buffer[562] ;
    input \data_buffer[563] ;
    input \data_buffer[564] ;
    input \data_buffer[568] ;
    input \data_buffer[160] ;
    input \data_buffer[569] ;
    input \data_buffer[570] ;
    input \data_buffer[571] ;
    input clk_c;
    input \data_buffer[572] ;
    input \data_buffer[576] ;
    input \data_buffer[577] ;
    input \data_buffer[416] ;
    input \data_buffer[578] ;
    input \data_buffer[579] ;
    input \data_buffer[580] ;
    input \data_buffer[584] ;
    input \data_buffer[585] ;
    input \data_buffer[586] ;
    input \data_buffer[587] ;
    input \data_buffer[588] ;
    input \data_buffer[592] ;
    input \data_buffer[593] ;
    input \data_buffer[594] ;
    input \data_buffer[595] ;
    input \data_buffer[596] ;
    input \data_buffer[600] ;
    input \data_buffer[601] ;
    input \data_buffer[602] ;
    input \data_buffer[603] ;
    input \data_buffer[604] ;
    input \data_buffer[608] ;
    input \data_buffer[609] ;
    input \data_buffer[610] ;
    input \data_buffer[611] ;
    input \data_buffer[612] ;
    input \data_buffer[616] ;
    input \data_buffer[617] ;
    input \data_buffer[618] ;
    input \data_buffer[619] ;
    input \data_buffer[620] ;
    input \data_buffer[624] ;
    input \data_buffer[625] ;
    input \data_buffer[626] ;
    input \data_buffer[627] ;
    input \data_buffer[628] ;
    output [9:0]data_length_reg;
    output n15;
    input \data_buffer[632] ;
    input \data_buffer[633] ;
    input \data_buffer[634] ;
    input \data_buffer[635] ;
    input \data_buffer[636] ;
    input \data_buffer[640] ;
    input \data_buffer[641] ;
    input \data_buffer[642] ;
    input \data_buffer[643] ;
    input \data_buffer[644] ;
    input \data_buffer[648] ;
    input \data_buffer[649] ;
    input \data_buffer[650] ;
    input \data_buffer[651] ;
    input \data_buffer[652] ;
    input \data_buffer[656] ;
    input \data_buffer[657] ;
    input \data_buffer[658] ;
    input \data_buffer[659] ;
    input \data_buffer[660] ;
    input \data_buffer[664] ;
    input \data_buffer[665] ;
    input \data_buffer[666] ;
    input \data_buffer[667] ;
    input \data_buffer[668] ;
    input \data_buffer[672] ;
    input \data_buffer[673] ;
    input \data_buffer[674] ;
    input \data_buffer[675] ;
    input \data_buffer[676] ;
    input \data_buffer[680] ;
    input \data_buffer[681] ;
    input \data_buffer[682] ;
    input \data_buffer[683] ;
    input \data_buffer[684] ;
    input \data_buffer[688] ;
    input \data_buffer[689] ;
    input \data_buffer[690] ;
    input \data_buffer[691] ;
    input \data_buffer[692] ;
    input \data_buffer[696] ;
    input \data_buffer[697] ;
    input \data_buffer[698] ;
    input \data_buffer[699] ;
    input \data_buffer[700] ;
    input \data_buffer[704] ;
    input \data_buffer[705] ;
    input \data_buffer[706] ;
    input \data_buffer[707] ;
    input \data_buffer[708] ;
    input \data_buffer[712] ;
    input \data_buffer[713] ;
    input \data_buffer[714] ;
    input \data_buffer[715] ;
    input \data_buffer[716] ;
    input \data_buffer[720] ;
    input \data_buffer[161] ;
    input \data_buffer[721] ;
    input \data_buffer[722] ;
    input \data_buffer[723] ;
    input \data_buffer[724] ;
    input \data_buffer[728] ;
    input \data_buffer[729] ;
    input \data_buffer[730] ;
    input \data_buffer[731] ;
    input \data_buffer[732] ;
    input \data_buffer[736] ;
    input \data_buffer[737] ;
    input \data_buffer[162] ;
    input \data_buffer[738] ;
    input \data_buffer[739] ;
    input \data_buffer[740] ;
    input \data_buffer[744] ;
    input \data_buffer[163] ;
    input \data_buffer[745] ;
    input \data_buffer[746] ;
    input \data_buffer[747] ;
    input \data_buffer[748] ;
    input \data_buffer[752] ;
    input \data_buffer[753] ;
    input \data_buffer[754] ;
    input \data_buffer[755] ;
    input \data_buffer[756] ;
    input \data_buffer[760] ;
    input \data_buffer[761] ;
    input \data_buffer[762] ;
    input \data_buffer[763] ;
    input \data_buffer[764] ;
    input \data_buffer[768] ;
    input \data_buffer[769] ;
    input \data_buffer[770] ;
    input \data_buffer[771] ;
    input \data_buffer[772] ;
    input \data_buffer[776] ;
    input \data_buffer[777] ;
    input \data_buffer[778] ;
    input \data_buffer[779] ;
    input \data_buffer[780] ;
    input \data_buffer[784] ;
    input \data_buffer[785] ;
    input \data_buffer[786] ;
    input \data_buffer[787] ;
    input \data_buffer[788] ;
    input \data_buffer[792] ;
    input \data_buffer[793] ;
    input \data_buffer[794] ;
    input \data_buffer[164] ;
    input \data_buffer[795] ;
    input \data_buffer[796] ;
    input \data_buffer[800] ;
    input \data_buffer[801] ;
    input \data_buffer[802] ;
    input \data_buffer[803] ;
    input \data_buffer[804] ;
    input \data_buffer[808] ;
    input \data_buffer[809] ;
    input \data_buffer[810] ;
    input \data_buffer[811] ;
    input \data_buffer[812] ;
    input \data_buffer[816] ;
    input \data_buffer[817] ;
    input \data_buffer[818] ;
    input \data_buffer[819] ;
    input \data_buffer[820] ;
    input \data_buffer[824] ;
    input \data_buffer[825] ;
    input \data_buffer[826] ;
    input \data_buffer[827] ;
    input \data_buffer[828] ;
    input \data_buffer[832] ;
    input \data_buffer[833] ;
    input \data_buffer[834] ;
    input \data_buffer[835] ;
    input \data_buffer[836] ;
    input \data_buffer[840] ;
    input \data_buffer[841] ;
    input \data_buffer[842] ;
    input \data_buffer[843] ;
    input \data_buffer[844] ;
    input \data_buffer[848] ;
    input \data_buffer[849] ;
    input \data_buffer[850] ;
    input \data_buffer[851] ;
    input \data_buffer[852] ;
    input \data_buffer[856] ;
    input \data_buffer[857] ;
    input \data_buffer[858] ;
    input \data_buffer[859] ;
    input \data_buffer[860] ;
    input \data_buffer[864] ;
    input \data_buffer[865] ;
    input \data_buffer[866] ;
    input \data_buffer[867] ;
    input \data_buffer[868] ;
    input \data_buffer[872] ;
    input \data_buffer[873] ;
    input \data_buffer[874] ;
    input \data_buffer[875] ;
    input \data_buffer[876] ;
    input \data_buffer[880] ;
    input \data_buffer[881] ;
    input \data_buffer[882] ;
    input \data_buffer[883] ;
    input \data_buffer[884] ;
    input \data_buffer[888] ;
    input \data_buffer[889] ;
    input \data_buffer[890] ;
    input \data_buffer[891] ;
    input \data_buffer[892] ;
    input \data_buffer[386] ;
    input \data_buffer[896] ;
    input \data_buffer[897] ;
    input \data_buffer[898] ;
    input \data_buffer[899] ;
    input \data_buffer[900] ;
    input \data_buffer[904] ;
    input \data_buffer[905] ;
    input \data_buffer[906] ;
    input \data_buffer[907] ;
    input \data_buffer[908] ;
    input \data_buffer[912] ;
    input \data_buffer[913] ;
    input \data_buffer[914] ;
    input \data_buffer[915] ;
    input \data_buffer[916] ;
    input \data_buffer[920] ;
    input \data_buffer[921] ;
    input \data_buffer[922] ;
    input \data_buffer[923] ;
    input \data_buffer[924] ;
    input \data_buffer[928] ;
    input \data_buffer[929] ;
    input \data_buffer[930] ;
    input \data_buffer[931] ;
    input \data_buffer[932] ;
    input \data_buffer[168] ;
    input \data_buffer[936] ;
    input \data_buffer[937] ;
    input \data_buffer[938] ;
    input \data_buffer[939] ;
    input \data_buffer[940] ;
    input \data_buffer[944] ;
    input \data_buffer[945] ;
    input \data_buffer[946] ;
    input \data_buffer[947] ;
    input \data_buffer[948] ;
    input \data_buffer[169] ;
    input \data_buffer[170] ;
    input \data_buffer[171] ;
    input \data_buffer[0] ;
    input \data_buffer[387] ;
    input \data_buffer[172] ;
    input \data_buffer[176] ;
    input \data_buffer[177] ;
    input \data_buffer[178] ;
    input \data_buffer[956] ;
    input \data_buffer[179] ;
    input \data_buffer[1] ;
    input \data_buffer[2] ;
    input \data_buffer[3] ;
    input \data_buffer[4] ;
    input \data_buffer[8] ;
    input \data_buffer[9] ;
    input \data_buffer[10] ;
    input \data_buffer[11] ;
    input \data_buffer[12] ;
    input \data_buffer[16] ;
    input \data_buffer[17] ;
    input \data_buffer[18] ;
    input \data_buffer[19] ;
    input \data_buffer[20] ;
    input \data_buffer[24] ;
    input \data_buffer[25] ;
    input \data_buffer[26] ;
    input \data_buffer[27] ;
    input \data_buffer[28] ;
    input \data_buffer[32] ;
    input \data_buffer[33] ;
    input \data_buffer[955] ;
    input \data_buffer[34] ;
    input \data_buffer[35] ;
    input \data_buffer[36] ;
    input \data_buffer[40] ;
    input \data_buffer[41] ;
    input \data_buffer[42] ;
    input \data_buffer[43] ;
    input \data_buffer[44] ;
    input \data_buffer[48] ;
    input \data_buffer[49] ;
    input \data_buffer[50] ;
    input \data_buffer[51] ;
    input \data_buffer[52] ;
    input \data_buffer[56] ;
    input \data_buffer[57] ;
    input \data_buffer[58] ;
    input \data_buffer[954] ;
    input \data_buffer[59] ;
    input \data_buffer[60] ;
    input \data_buffer[388] ;
    input \data_buffer[64] ;
    input \data_buffer[953] ;
    input \data_buffer[952] ;
    input \data_buffer[65] ;
    input \data_buffer[180] ;
    input \data_buffer[66] ;
    input \data_buffer[67] ;
    input \data_buffer[68] ;
    input \data_buffer[72] ;
    input \data_buffer[73] ;
    input \data_buffer[74] ;
    input \data_buffer[75] ;
    input \data_buffer[76] ;
    input \data_buffer[80] ;
    input \data_buffer[81] ;
    input \data_buffer[82] ;
    input \data_buffer[83] ;
    input \data_buffer[84] ;
    input \data_buffer[88] ;
    input \data_buffer[184] ;
    input \data_buffer[89] ;
    input \data_buffer[90] ;
    input \data_buffer[185] ;
    input \data_buffer[91] ;
    input \data_buffer[92] ;
    input \data_buffer[96] ;
    input \data_buffer[97] ;
    input \data_buffer[98] ;
    input \data_buffer[99] ;
    input \data_buffer[100] ;
    input \data_buffer[186] ;
    input \data_buffer[104] ;
    input \data_buffer[105] ;
    input \data_buffer[106] ;
    input \data_buffer[107] ;
    input \data_buffer[108] ;
    input \data_buffer[112] ;
    input \data_buffer[113] ;
    input \data_buffer[114] ;
    input \data_buffer[115] ;
    input \data_buffer[116] ;
    input \data_buffer[120] ;
    input \data_buffer[121] ;
    input \data_buffer[122] ;
    input \data_buffer[123] ;
    input \data_buffer[124] ;
    input \data_buffer[128] ;
    input \data_buffer[129] ;
    input \data_buffer[187] ;
    input \data_buffer[130] ;
    input \data_buffer[131] ;
    input \data_buffer[132] ;
    input \data_buffer[136] ;
    input \data_buffer[137] ;
    input \data_buffer[138] ;
    input \data_buffer[139] ;
    input \data_buffer[140] ;
    input \data_buffer[144] ;
    input \data_buffer[145] ;
    input \data_buffer[146] ;
    input \data_buffer[147] ;
    input \data_buffer[148] ;
    input \data_buffer[152] ;
    input \data_buffer[153] ;
    input \data_buffer[154] ;
    input \data_buffer[155] ;
    input \data_buffer[156] ;
    input \data_buffer[188] ;
    input \data_buffer[392] ;
    input \data_buffer[393] ;
    input \data_buffer[394] ;
    input \data_buffer[192] ;
    input \data_buffer[193] ;
    input \data_buffer[194] ;
    input \data_buffer[195] ;
    input \data_buffer[196] ;
    input \data_buffer[200] ;
    input \data_buffer[395] ;
    input \data_buffer[396] ;
    input \data_buffer[201] ;
    input \data_buffer[202] ;
    input \data_buffer[203] ;
    input \data_buffer[204] ;
    input \data_buffer[208] ;
    input \data_buffer[417] ;
    input \data_buffer[418] ;
    input \data_buffer[419] ;
    input \data_buffer[420] ;
    input \data_buffer[400] ;
    input \data_buffer[401] ;
    input \data_buffer[209] ;
    input \data_buffer[210] ;
    input \data_buffer[424] ;
    input \data_buffer[211] ;
    input \data_buffer[425] ;
    input \data_buffer[212] ;
    input \data_buffer[426] ;
    input \data_buffer[402] ;
    input \data_buffer[427] ;
    input \data_buffer[428] ;
    input \data_buffer[216] ;
    input \data_buffer[217] ;
    input \data_buffer[218] ;
    input \data_buffer[219] ;
    input \data_buffer[432] ;
    input \data_buffer[433] ;
    input \data_buffer[220] ;
    input \data_buffer[434] ;
    input \data_buffer[435] ;
    input \data_buffer[436] ;
    input \data_buffer[440] ;
    input \data_buffer[224] ;
    input \data_buffer[225] ;
    input \data_buffer[441] ;
    input \data_buffer[403] ;
    input \data_buffer[226] ;
    input \data_buffer[227] ;
    input \data_buffer[228] ;
    input \data_buffer[232] ;
    input \data_buffer[233] ;
    input \data_buffer[234] ;
    input \data_buffer[442] ;
    input \data_buffer[443] ;
    input \data_buffer[404] ;
    input \data_buffer[444] ;
    input \data_buffer[235] ;
    input \data_buffer[236] ;
    input \data_buffer[408] ;
    input \data_buffer[240] ;
    input \data_buffer[409] ;
    input \data_buffer[241] ;
    input \data_buffer[448] ;
    input \data_buffer[242] ;
    input \data_buffer[449] ;
    input \data_buffer[450] ;
    input \data_buffer[243] ;
    input \data_buffer[451] ;
    input \data_buffer[244] ;
    input \data_buffer[248] ;
    input \data_buffer[452] ;
    input \data_buffer[249] ;
    input \data_buffer[250] ;
    input \data_buffer[251] ;
    input \data_buffer[252] ;
    input \data_buffer[256] ;
    input \data_buffer[257] ;
    input \data_buffer[258] ;
    input \data_buffer[259] ;
    input \data_buffer[260] ;
    input \data_buffer[264] ;
    input \data_buffer[265] ;
    input \data_buffer[266] ;
    input \data_buffer[267] ;
    input \data_buffer[268] ;
    input \data_buffer[272] ;
    input \data_buffer[456] ;
    input \data_buffer[273] ;
    input \data_buffer[274] ;
    input \data_buffer[457] ;
    input \data_buffer[275] ;
    input \data_buffer[276] ;
    input \data_buffer[458] ;
    input [9:0]data_length;
    input GND_net;
    input \data_buffer[280] ;
    input \data_buffer[459] ;
    input \data_buffer[460] ;
    input \data_buffer[281] ;
    input \data_buffer[282] ;
    input \data_buffer[283] ;
    input \data_buffer[284] ;
    input \data_buffer[288] ;
    input \data_buffer[464] ;
    input \data_buffer[289] ;
    input \data_buffer[465] ;
    input \data_buffer[290] ;
    input \data_buffer[466] ;
    input \data_buffer[291] ;
    input \data_buffer[292] ;
    input \data_buffer[296] ;
    input \data_buffer[467] ;
    input \data_buffer[297] ;
    input \data_buffer[298] ;
    input \data_buffer[468] ;
    input \data_buffer[472] ;
    input \data_buffer[299] ;
    input \data_buffer[300] ;
    input \data_buffer[304] ;
    input \data_buffer[305] ;
    input \data_buffer[306] ;
    input \data_buffer[307] ;
    input \data_buffer[308] ;
    input \data_buffer[312] ;
    input \data_buffer[473] ;
    input \data_buffer[313] ;
    input \data_buffer[314] ;
    input \data_buffer[315] ;
    input \data_buffer[474] ;
    input \data_buffer[316] ;
    input \data_buffer[475] ;
    input \data_buffer[320] ;
    input \data_buffer[321] ;
    input \data_buffer[476] ;
    input \data_buffer[480] ;
    input \data_buffer[322] ;
    input \data_buffer[323] ;
    input \data_buffer[324] ;
    input \data_buffer[481] ;
    input \data_buffer[328] ;
    input \data_buffer[329] ;
    input \data_buffer[330] ;
    input \data_buffer[331] ;
    input \data_buffer[482] ;
    input \data_buffer[483] ;
    input \data_buffer[484] ;
    input \data_buffer[332] ;
    input \data_buffer[488] ;
    input \data_buffer[336] ;
    input \data_buffer[337] ;
    input \data_buffer[489] ;
    input \data_buffer[338] ;
    input \data_buffer[490] ;
    input \data_buffer[339] ;
    input \data_buffer[491] ;
    input \data_buffer[340] ;
    input \data_buffer[344] ;
    input \data_buffer[492] ;
    input \data_buffer[345] ;
    input \data_buffer[496] ;
    input \data_buffer[497] ;
    input \data_buffer[346] ;
    input \data_buffer[347] ;
    input \data_buffer[498] ;
    input \data_buffer[499] ;
    input \data_buffer[500] ;
    input \data_buffer[348] ;
    input \data_buffer[352] ;
    input \data_buffer[353] ;
    input \data_buffer[354] ;
    input \data_buffer[355] ;
    input \data_buffer[356] ;
    input \data_buffer[504] ;
    input \data_buffer[360] ;
    input \data_buffer[361] ;
    input \data_buffer[505] ;
    input \data_buffer[506] ;
    input \data_buffer[362] ;
    input \data_buffer[507] ;
    input \data_buffer[363] ;
    input \data_buffer[508] ;
    input \data_buffer[364] ;
    input \data_buffer[368] ;
    input \data_buffer[369] ;
    input \data_buffer[512] ;
    input \data_buffer[513] ;
    input \data_buffer[514] ;
    input \data_buffer[515] ;
    input \data_buffer[370] ;
    input \data_buffer[516] ;
    input \data_buffer[520] ;
    input \data_buffer[371] ;
    input \data_buffer[521] ;
    input \data_buffer[372] ;
    input \data_buffer[522] ;
    input \data_buffer[523] ;
    input \data_buffer[524] ;
    input \data_buffer[376] ;
    input \data_buffer[528] ;
    input \data_buffer[529] ;
    input \data_buffer[530] ;
    input \data_buffer[531] ;
    input \data_buffer[532] ;
    input \data_buffer[536] ;
    input \data_buffer[537] ;
    input \data_buffer[377] ;
    input \data_buffer[378] ;
    input \data_buffer[379] ;
    input \data_buffer[380] ;
    input \data_buffer[410] ;
    input \data_buffer[411] ;
    input \data_buffer[412] ;
    input \data_buffer[384] ;
    input \data_buffer[385] ;
    output piano_out_c;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // g:/fpga/mxo2/system/project/system_top.v(2[15:18])
    wire [959:0]data_buffer_reg;   // g:/fpga/mxo2/system/project/beeper_control.v(31[23:38])
    wire [959:0]data_buffer_reg_959__N_3020;
    
    wire clk_c_enable_799, n25588;
    wire [23:0]cnt;   // g:/fpga/mxo2/system/project/beeper_control.v(12[14:17])
    wire [23:0]n101;
    wire [9:0]n45;
    
    wire clk_c_enable_899, clk_c_enable_950, clk_c_enable_1000, clk_c_enable_1200, 
        clk_c_enable_849, clk_c_enable_1050, clk_c_enable_1100, clk_c_enable_1150, 
        clk_c_enable_1250, clk_c_enable_1304, clk_c_enable_1414, n15_adj_5036;
    wire [9:0]data_length_reg_c;   // g:/fpga/mxo2/system/project/beeper_control.v(22[21:36])
    
    wire n14, n23729, n21027, n24165, n23723, n23809, n17, n16, 
        n25623, n12089, n3057, n2025, n20546, n20545, n20544, 
        n20543, n20542, n25562, n20538, n20537, n20536, n20535, 
        n20534, n20533, n20532, n20531, n20530, n20529, n20528, 
        n20527;
    
    LUT4 data_buffer_reg_959__I_0_i539_3_lut (.A(data_buffer_reg[546]), .B(\data_buffer[538] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[538])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i539_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i540_3_lut (.A(data_buffer_reg[547]), .B(\data_buffer[539] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[539])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i540_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i541_3_lut (.A(data_buffer_reg[548]), .B(\data_buffer[540] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[540])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i541_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i545_3_lut (.A(data_buffer_reg[552]), .B(\data_buffer[544] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[544])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i545_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i546_3_lut (.A(data_buffer_reg[553]), .B(\data_buffer[545] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[545])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i546_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i547_3_lut (.A(data_buffer_reg[554]), .B(\data_buffer[546] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[546])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i547_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i548_3_lut (.A(data_buffer_reg[555]), .B(\data_buffer[547] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[547])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i548_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i549_3_lut (.A(data_buffer_reg[556]), .B(\data_buffer[548] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[548])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i549_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i553_3_lut (.A(data_buffer_reg[560]), .B(\data_buffer[552] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[552])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i553_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i554_3_lut (.A(data_buffer_reg[561]), .B(\data_buffer[553] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[553])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i554_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i555_3_lut (.A(data_buffer_reg[562]), .B(\data_buffer[554] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[554])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i555_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i556_3_lut (.A(data_buffer_reg[563]), .B(\data_buffer[555] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[555])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i556_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i557_3_lut (.A(data_buffer_reg[564]), .B(\data_buffer[556] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[556])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i557_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i561_3_lut (.A(data_buffer_reg[568]), .B(\data_buffer[560] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[560])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i561_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i562_3_lut (.A(data_buffer_reg[569]), .B(\data_buffer[561] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[561])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i562_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i563_3_lut (.A(data_buffer_reg[570]), .B(\data_buffer[562] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[562])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i563_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i564_3_lut (.A(data_buffer_reg[571]), .B(\data_buffer[563] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[563])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i564_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i565_3_lut (.A(data_buffer_reg[572]), .B(\data_buffer[564] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[564])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i565_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i569_3_lut (.A(data_buffer_reg[576]), .B(\data_buffer[568] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[568])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i569_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i161_3_lut (.A(data_buffer_reg[168]), .B(\data_buffer[160] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[160])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i161_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i570_3_lut (.A(data_buffer_reg[577]), .B(\data_buffer[569] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[569])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i570_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i571_3_lut (.A(data_buffer_reg[578]), .B(\data_buffer[570] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[570])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i571_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i572_3_lut (.A(data_buffer_reg[579]), .B(\data_buffer[571] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[571])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i572_3_lut.init = 16'hcaca;
    FD1P3AX data_buffer_reg_i0 (.D(data_buffer_reg_959__N_3020[0]), .SP(clk_c_enable_799), 
            .CK(clk_c), .Q(data_buffer_reg[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i0.GSR = "ENABLED";
    LUT4 data_buffer_reg_959__I_0_i573_3_lut (.A(data_buffer_reg[580]), .B(\data_buffer[572] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[572])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i573_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i577_3_lut (.A(data_buffer_reg[584]), .B(\data_buffer[576] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[576])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i577_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i578_3_lut (.A(data_buffer_reg[585]), .B(\data_buffer[577] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[577])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i578_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i417_3_lut (.A(data_buffer_reg[424]), .B(\data_buffer[416] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[416])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i417_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i579_3_lut (.A(data_buffer_reg[586]), .B(\data_buffer[578] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[578])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i579_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i580_3_lut (.A(data_buffer_reg[587]), .B(\data_buffer[579] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[579])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i580_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i581_3_lut (.A(data_buffer_reg[588]), .B(\data_buffer[580] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[580])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i581_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i585_3_lut (.A(data_buffer_reg[592]), .B(\data_buffer[584] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[584])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i585_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i586_3_lut (.A(data_buffer_reg[593]), .B(\data_buffer[585] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[585])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i586_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i587_3_lut (.A(data_buffer_reg[594]), .B(\data_buffer[586] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[586])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i587_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i588_3_lut (.A(data_buffer_reg[595]), .B(\data_buffer[587] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[587])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i588_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i589_3_lut (.A(data_buffer_reg[596]), .B(\data_buffer[588] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[588])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i589_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i593_3_lut (.A(data_buffer_reg[600]), .B(\data_buffer[592] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[592])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i593_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i594_3_lut (.A(data_buffer_reg[601]), .B(\data_buffer[593] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[593])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i594_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i595_3_lut (.A(data_buffer_reg[602]), .B(\data_buffer[594] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[594])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i595_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i596_3_lut (.A(data_buffer_reg[603]), .B(\data_buffer[595] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[595])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i596_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i597_3_lut (.A(data_buffer_reg[604]), .B(\data_buffer[596] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[596])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i597_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i601_3_lut (.A(data_buffer_reg[608]), .B(\data_buffer[600] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[600])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i601_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i602_3_lut (.A(data_buffer_reg[609]), .B(\data_buffer[601] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[601])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i602_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i603_3_lut (.A(data_buffer_reg[610]), .B(\data_buffer[602] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[602])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i603_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i604_3_lut (.A(data_buffer_reg[611]), .B(\data_buffer[603] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[603])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i604_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i605_3_lut (.A(data_buffer_reg[612]), .B(\data_buffer[604] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[604])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i605_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i609_3_lut (.A(data_buffer_reg[616]), .B(\data_buffer[608] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[608])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i609_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i610_3_lut (.A(data_buffer_reg[617]), .B(\data_buffer[609] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[609])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i610_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i611_3_lut (.A(data_buffer_reg[618]), .B(\data_buffer[610] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[610])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i611_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i612_3_lut (.A(data_buffer_reg[619]), .B(\data_buffer[611] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[611])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i612_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i613_3_lut (.A(data_buffer_reg[620]), .B(\data_buffer[612] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[612])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i613_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i617_3_lut (.A(data_buffer_reg[624]), .B(\data_buffer[616] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[616])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i617_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i618_3_lut (.A(data_buffer_reg[625]), .B(\data_buffer[617] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[617])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i618_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i619_3_lut (.A(data_buffer_reg[626]), .B(\data_buffer[618] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[618])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i619_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i620_3_lut (.A(data_buffer_reg[627]), .B(\data_buffer[619] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[619])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i620_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i621_3_lut (.A(data_buffer_reg[628]), .B(\data_buffer[620] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[620])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i621_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i625_3_lut (.A(data_buffer_reg[632]), .B(\data_buffer[624] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[624])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i625_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i626_3_lut (.A(data_buffer_reg[633]), .B(\data_buffer[625] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[625])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i626_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i627_3_lut (.A(data_buffer_reg[634]), .B(\data_buffer[626] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[626])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i627_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i628_3_lut (.A(data_buffer_reg[635]), .B(\data_buffer[627] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[627])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i628_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i629_3_lut (.A(data_buffer_reg[636]), .B(\data_buffer[628] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[628])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i629_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_3_lut_4_lut_rep_485 (.A(data_length_reg[0]), .B(n15), 
         .C(n26793), .D(n25588), .Z(clk_c_enable_799)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i1_2_lut_3_lut_3_lut_4_lut_rep_485.init = 16'hfef0;
    LUT4 data_buffer_reg_959__I_0_i633_3_lut (.A(data_buffer_reg[640]), .B(\data_buffer[632] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[632])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i633_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i634_3_lut (.A(data_buffer_reg[641]), .B(\data_buffer[633] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[633])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i634_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i635_3_lut (.A(data_buffer_reg[642]), .B(\data_buffer[634] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[634])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i635_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i636_3_lut (.A(data_buffer_reg[643]), .B(\data_buffer[635] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[635])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i636_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i637_3_lut (.A(data_buffer_reg[644]), .B(\data_buffer[636] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[636])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i637_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i641_3_lut (.A(data_buffer_reg[648]), .B(\data_buffer[640] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[640])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i641_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i642_3_lut (.A(data_buffer_reg[649]), .B(\data_buffer[641] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[641])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i642_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i643_3_lut (.A(data_buffer_reg[650]), .B(\data_buffer[642] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[642])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i643_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i644_3_lut (.A(data_buffer_reg[651]), .B(\data_buffer[643] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[643])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i644_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i645_3_lut (.A(data_buffer_reg[652]), .B(\data_buffer[644] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[644])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i645_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i649_3_lut (.A(data_buffer_reg[656]), .B(\data_buffer[648] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[648])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i649_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i650_3_lut (.A(data_buffer_reg[657]), .B(\data_buffer[649] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[649])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i650_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i651_3_lut (.A(data_buffer_reg[658]), .B(\data_buffer[650] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[650])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i651_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i652_3_lut (.A(data_buffer_reg[659]), .B(\data_buffer[651] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[651])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i652_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i653_3_lut (.A(data_buffer_reg[660]), .B(\data_buffer[652] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[652])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i653_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i657_3_lut (.A(data_buffer_reg[664]), .B(\data_buffer[656] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[656])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i657_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i658_3_lut (.A(data_buffer_reg[665]), .B(\data_buffer[657] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[657])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i658_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i659_3_lut (.A(data_buffer_reg[666]), .B(\data_buffer[658] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[658])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i659_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i660_3_lut (.A(data_buffer_reg[667]), .B(\data_buffer[659] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[659])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i660_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i661_3_lut (.A(data_buffer_reg[668]), .B(\data_buffer[660] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[660])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i661_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i665_3_lut (.A(data_buffer_reg[672]), .B(\data_buffer[664] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[664])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i665_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i666_3_lut (.A(data_buffer_reg[673]), .B(\data_buffer[665] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[665])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i666_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i667_3_lut (.A(data_buffer_reg[674]), .B(\data_buffer[666] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[666])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i667_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i668_3_lut (.A(data_buffer_reg[675]), .B(\data_buffer[667] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[667])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i668_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i669_3_lut (.A(data_buffer_reg[676]), .B(\data_buffer[668] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[668])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i669_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i673_3_lut (.A(data_buffer_reg[680]), .B(\data_buffer[672] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[672])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i673_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i674_3_lut (.A(data_buffer_reg[681]), .B(\data_buffer[673] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[673])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i674_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i675_3_lut (.A(data_buffer_reg[682]), .B(\data_buffer[674] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[674])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i675_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i676_3_lut (.A(data_buffer_reg[683]), .B(\data_buffer[675] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[675])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i676_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i677_3_lut (.A(data_buffer_reg[684]), .B(\data_buffer[676] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[676])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i677_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i681_3_lut (.A(data_buffer_reg[688]), .B(\data_buffer[680] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[680])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i681_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i682_3_lut (.A(data_buffer_reg[689]), .B(\data_buffer[681] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[681])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i682_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i683_3_lut (.A(data_buffer_reg[690]), .B(\data_buffer[682] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[682])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i683_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i684_3_lut (.A(data_buffer_reg[691]), .B(\data_buffer[683] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[683])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i684_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i685_3_lut (.A(data_buffer_reg[692]), .B(\data_buffer[684] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[684])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i685_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i689_3_lut (.A(data_buffer_reg[696]), .B(\data_buffer[688] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[688])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i689_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i690_3_lut (.A(data_buffer_reg[697]), .B(\data_buffer[689] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[689])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i690_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i691_3_lut (.A(data_buffer_reg[698]), .B(\data_buffer[690] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[690])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i691_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i692_3_lut (.A(data_buffer_reg[699]), .B(\data_buffer[691] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[691])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i692_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i693_3_lut (.A(data_buffer_reg[700]), .B(\data_buffer[692] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[692])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i693_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i697_3_lut (.A(data_buffer_reg[704]), .B(\data_buffer[696] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[696])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i697_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i698_3_lut (.A(data_buffer_reg[705]), .B(\data_buffer[697] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[697])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i698_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i699_3_lut (.A(data_buffer_reg[706]), .B(\data_buffer[698] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[698])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i699_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i700_3_lut (.A(data_buffer_reg[707]), .B(\data_buffer[699] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[699])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i700_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i701_3_lut (.A(data_buffer_reg[708]), .B(\data_buffer[700] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[700])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i701_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i705_3_lut (.A(data_buffer_reg[712]), .B(\data_buffer[704] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[704])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i705_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i706_3_lut (.A(data_buffer_reg[713]), .B(\data_buffer[705] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[705])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i706_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i707_3_lut (.A(data_buffer_reg[714]), .B(\data_buffer[706] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[706])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i707_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i708_3_lut (.A(data_buffer_reg[715]), .B(\data_buffer[707] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[707])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i708_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i709_3_lut (.A(data_buffer_reg[716]), .B(\data_buffer[708] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[708])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i709_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i713_3_lut (.A(data_buffer_reg[720]), .B(\data_buffer[712] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[712])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i713_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i714_3_lut (.A(data_buffer_reg[721]), .B(\data_buffer[713] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[713])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i714_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i715_3_lut (.A(data_buffer_reg[722]), .B(\data_buffer[714] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[714])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i715_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i716_3_lut (.A(data_buffer_reg[723]), .B(\data_buffer[715] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[715])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i716_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i717_3_lut (.A(data_buffer_reg[724]), .B(\data_buffer[716] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[716])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i717_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i721_3_lut (.A(data_buffer_reg[728]), .B(\data_buffer[720] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[720])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i721_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i162_3_lut (.A(data_buffer_reg[169]), .B(\data_buffer[161] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[161])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i162_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i722_3_lut (.A(data_buffer_reg[729]), .B(\data_buffer[721] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[721])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i722_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i723_3_lut (.A(data_buffer_reg[730]), .B(\data_buffer[722] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[722])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i723_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i724_3_lut (.A(data_buffer_reg[731]), .B(\data_buffer[723] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[723])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i724_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i725_3_lut (.A(data_buffer_reg[732]), .B(\data_buffer[724] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[724])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i725_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i729_3_lut (.A(data_buffer_reg[736]), .B(\data_buffer[728] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[728])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i729_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i730_3_lut (.A(data_buffer_reg[737]), .B(\data_buffer[729] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[729])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i730_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i731_3_lut (.A(data_buffer_reg[738]), .B(\data_buffer[730] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[730])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i731_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i732_3_lut (.A(data_buffer_reg[739]), .B(\data_buffer[731] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[731])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i732_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i733_3_lut (.A(data_buffer_reg[740]), .B(\data_buffer[732] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[732])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i733_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i737_3_lut (.A(data_buffer_reg[744]), .B(\data_buffer[736] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[736])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i737_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i738_3_lut (.A(data_buffer_reg[745]), .B(\data_buffer[737] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[737])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i738_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i163_3_lut (.A(data_buffer_reg[170]), .B(\data_buffer[162] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[162])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i163_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i739_3_lut (.A(data_buffer_reg[746]), .B(\data_buffer[738] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[738])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i739_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i740_3_lut (.A(data_buffer_reg[747]), .B(\data_buffer[739] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[739])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i740_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i741_3_lut (.A(data_buffer_reg[748]), .B(\data_buffer[740] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[740])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i741_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i745_3_lut (.A(data_buffer_reg[752]), .B(\data_buffer[744] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[744])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i745_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i164_3_lut (.A(data_buffer_reg[171]), .B(\data_buffer[163] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[163])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i164_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i746_3_lut (.A(data_buffer_reg[753]), .B(\data_buffer[745] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[745])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i746_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i747_3_lut (.A(data_buffer_reg[754]), .B(\data_buffer[746] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[746])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i747_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i748_3_lut (.A(data_buffer_reg[755]), .B(\data_buffer[747] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[747])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i748_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i749_3_lut (.A(data_buffer_reg[756]), .B(\data_buffer[748] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[748])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i749_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i753_3_lut (.A(data_buffer_reg[760]), .B(\data_buffer[752] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[752])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i753_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i754_3_lut (.A(data_buffer_reg[761]), .B(\data_buffer[753] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[753])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i754_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i755_3_lut (.A(data_buffer_reg[762]), .B(\data_buffer[754] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[754])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i755_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i756_3_lut (.A(data_buffer_reg[763]), .B(\data_buffer[755] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[755])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i756_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i757_3_lut (.A(data_buffer_reg[764]), .B(\data_buffer[756] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[756])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i757_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i761_3_lut (.A(data_buffer_reg[768]), .B(\data_buffer[760] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[760])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i761_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i762_3_lut (.A(data_buffer_reg[769]), .B(\data_buffer[761] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[761])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i762_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i763_3_lut (.A(data_buffer_reg[770]), .B(\data_buffer[762] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[762])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i763_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i764_3_lut (.A(data_buffer_reg[771]), .B(\data_buffer[763] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[763])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i764_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i765_3_lut (.A(data_buffer_reg[772]), .B(\data_buffer[764] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[764])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i765_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i769_3_lut (.A(data_buffer_reg[776]), .B(\data_buffer[768] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[768])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i769_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i770_3_lut (.A(data_buffer_reg[777]), .B(\data_buffer[769] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[769])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i770_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i771_3_lut (.A(data_buffer_reg[778]), .B(\data_buffer[770] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[770])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i771_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i772_3_lut (.A(data_buffer_reg[779]), .B(\data_buffer[771] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[771])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i772_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i773_3_lut (.A(data_buffer_reg[780]), .B(\data_buffer[772] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[772])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i773_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i777_3_lut (.A(data_buffer_reg[784]), .B(\data_buffer[776] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[776])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i777_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i778_3_lut (.A(data_buffer_reg[785]), .B(\data_buffer[777] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[777])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i778_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i779_3_lut (.A(data_buffer_reg[786]), .B(\data_buffer[778] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[778])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i779_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i780_3_lut (.A(data_buffer_reg[787]), .B(\data_buffer[779] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[779])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i780_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i781_3_lut (.A(data_buffer_reg[788]), .B(\data_buffer[780] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[780])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i781_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i785_3_lut (.A(data_buffer_reg[792]), .B(\data_buffer[784] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[784])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i785_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i786_3_lut (.A(data_buffer_reg[793]), .B(\data_buffer[785] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[785])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i786_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i787_3_lut (.A(data_buffer_reg[794]), .B(\data_buffer[786] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[786])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i787_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i788_3_lut (.A(data_buffer_reg[795]), .B(\data_buffer[787] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[787])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i788_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i789_3_lut (.A(data_buffer_reg[796]), .B(\data_buffer[788] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[788])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i789_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i793_3_lut (.A(data_buffer_reg[800]), .B(\data_buffer[792] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[792])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i793_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i794_3_lut (.A(data_buffer_reg[801]), .B(\data_buffer[793] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[793])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i794_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i795_3_lut (.A(data_buffer_reg[802]), .B(\data_buffer[794] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[794])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i795_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i165_3_lut (.A(data_buffer_reg[172]), .B(\data_buffer[164] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[164])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i165_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i796_3_lut (.A(data_buffer_reg[803]), .B(\data_buffer[795] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[795])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i796_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i797_3_lut (.A(data_buffer_reg[804]), .B(\data_buffer[796] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[796])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i797_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i801_3_lut (.A(data_buffer_reg[808]), .B(\data_buffer[800] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[800])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i801_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i802_3_lut (.A(data_buffer_reg[809]), .B(\data_buffer[801] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[801])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i802_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i803_3_lut (.A(data_buffer_reg[810]), .B(\data_buffer[802] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[802])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i803_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i804_3_lut (.A(data_buffer_reg[811]), .B(\data_buffer[803] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[803])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i804_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i805_3_lut (.A(data_buffer_reg[812]), .B(\data_buffer[804] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[804])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i805_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i809_3_lut (.A(data_buffer_reg[816]), .B(\data_buffer[808] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[808])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i809_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i810_3_lut (.A(data_buffer_reg[817]), .B(\data_buffer[809] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[809])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i810_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i811_3_lut (.A(data_buffer_reg[818]), .B(\data_buffer[810] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[810])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i811_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i812_3_lut (.A(data_buffer_reg[819]), .B(\data_buffer[811] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[811])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i812_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i813_3_lut (.A(data_buffer_reg[820]), .B(\data_buffer[812] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[812])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i813_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i817_3_lut (.A(data_buffer_reg[824]), .B(\data_buffer[816] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[816])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i817_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i818_3_lut (.A(data_buffer_reg[825]), .B(\data_buffer[817] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[817])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i818_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i819_3_lut (.A(data_buffer_reg[826]), .B(\data_buffer[818] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[818])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i819_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i820_3_lut (.A(data_buffer_reg[827]), .B(\data_buffer[819] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[819])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i820_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i821_3_lut (.A(data_buffer_reg[828]), .B(\data_buffer[820] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[820])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i821_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i825_3_lut (.A(data_buffer_reg[832]), .B(\data_buffer[824] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[824])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i825_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i826_3_lut (.A(data_buffer_reg[833]), .B(\data_buffer[825] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[825])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i826_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i827_3_lut (.A(data_buffer_reg[834]), .B(\data_buffer[826] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[826])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i827_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i828_3_lut (.A(data_buffer_reg[835]), .B(\data_buffer[827] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[827])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i828_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i829_3_lut (.A(data_buffer_reg[836]), .B(\data_buffer[828] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[828])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i829_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i833_3_lut (.A(data_buffer_reg[840]), .B(\data_buffer[832] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[832])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i833_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i834_3_lut (.A(data_buffer_reg[841]), .B(\data_buffer[833] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[833])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i834_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i835_3_lut (.A(data_buffer_reg[842]), .B(\data_buffer[834] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[834])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i835_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i836_3_lut (.A(data_buffer_reg[843]), .B(\data_buffer[835] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[835])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i836_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i837_3_lut (.A(data_buffer_reg[844]), .B(\data_buffer[836] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[836])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i837_3_lut.init = 16'hcaca;
    FD1S3IX cnt_1981__i0 (.D(n101[0]), .CK(clk_c), .CD(n25588), .Q(cnt[0])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(19[16:26])
    defparam cnt_1981__i0.GSR = "ENABLED";
    LUT4 data_buffer_reg_959__I_0_i841_3_lut (.A(data_buffer_reg[848]), .B(\data_buffer[840] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[840])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i841_3_lut.init = 16'hcaca;
    FD1S3AX data_length_reg_1982__i0 (.D(n45[0]), .CK(clk_c), .Q(data_length_reg[0])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(29[28:50])
    defparam data_length_reg_1982__i0.GSR = "ENABLED";
    LUT4 data_buffer_reg_959__I_0_i842_3_lut (.A(data_buffer_reg[849]), .B(\data_buffer[841] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[841])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i842_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i843_3_lut (.A(data_buffer_reg[850]), .B(\data_buffer[842] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[842])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i843_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i844_3_lut (.A(data_buffer_reg[851]), .B(\data_buffer[843] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[843])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i844_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i845_3_lut (.A(data_buffer_reg[852]), .B(\data_buffer[844] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[844])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i845_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i849_3_lut (.A(data_buffer_reg[856]), .B(\data_buffer[848] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[848])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i849_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i850_3_lut (.A(data_buffer_reg[857]), .B(\data_buffer[849] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[849])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i850_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i851_3_lut (.A(data_buffer_reg[858]), .B(\data_buffer[850] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[850])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i851_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i852_3_lut (.A(data_buffer_reg[859]), .B(\data_buffer[851] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[851])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i852_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i853_3_lut (.A(data_buffer_reg[860]), .B(\data_buffer[852] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[852])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i853_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i857_3_lut (.A(data_buffer_reg[864]), .B(\data_buffer[856] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[856])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i857_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i858_3_lut (.A(data_buffer_reg[865]), .B(\data_buffer[857] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[857])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i858_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i859_3_lut (.A(data_buffer_reg[866]), .B(\data_buffer[858] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[858])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i859_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i860_3_lut (.A(data_buffer_reg[867]), .B(\data_buffer[859] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[859])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i860_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i861_3_lut (.A(data_buffer_reg[868]), .B(\data_buffer[860] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[860])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i861_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i865_3_lut (.A(data_buffer_reg[872]), .B(\data_buffer[864] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[864])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i865_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i866_3_lut (.A(data_buffer_reg[873]), .B(\data_buffer[865] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[865])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i866_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i867_3_lut (.A(data_buffer_reg[874]), .B(\data_buffer[866] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[866])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i867_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i868_3_lut (.A(data_buffer_reg[875]), .B(\data_buffer[867] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[867])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i868_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i869_3_lut (.A(data_buffer_reg[876]), .B(\data_buffer[868] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[868])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i869_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i873_3_lut (.A(data_buffer_reg[880]), .B(\data_buffer[872] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[872])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i873_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i874_3_lut (.A(data_buffer_reg[881]), .B(\data_buffer[873] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[873])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i874_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i875_3_lut (.A(data_buffer_reg[882]), .B(\data_buffer[874] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[874])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i875_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i876_3_lut (.A(data_buffer_reg[883]), .B(\data_buffer[875] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[875])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i876_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i877_3_lut (.A(data_buffer_reg[884]), .B(\data_buffer[876] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[876])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i877_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i881_3_lut (.A(data_buffer_reg[888]), .B(\data_buffer[880] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[880])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i881_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i882_3_lut (.A(data_buffer_reg[889]), .B(\data_buffer[881] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[881])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i882_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i883_3_lut (.A(data_buffer_reg[890]), .B(\data_buffer[882] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[882])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i883_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i884_3_lut (.A(data_buffer_reg[891]), .B(\data_buffer[883] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[883])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i884_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i885_3_lut (.A(data_buffer_reg[892]), .B(\data_buffer[884] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[884])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i885_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i889_3_lut (.A(data_buffer_reg[896]), .B(\data_buffer[888] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[888])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i889_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i890_3_lut (.A(data_buffer_reg[897]), .B(\data_buffer[889] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[889])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i890_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i891_3_lut (.A(data_buffer_reg[898]), .B(\data_buffer[890] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[890])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i891_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i892_3_lut (.A(data_buffer_reg[899]), .B(\data_buffer[891] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[891])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i892_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i893_3_lut (.A(data_buffer_reg[900]), .B(\data_buffer[892] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[892])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i893_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i387_3_lut (.A(data_buffer_reg[394]), .B(\data_buffer[386] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[386])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i387_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_3_lut_4_lut_rep_487 (.A(data_length_reg[0]), .B(n15), 
         .C(n26793), .D(n25588), .Z(clk_c_enable_899)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i1_2_lut_3_lut_3_lut_4_lut_rep_487.init = 16'hfef0;
    LUT4 data_buffer_reg_959__I_0_i897_3_lut (.A(data_buffer_reg[904]), .B(\data_buffer[896] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[896])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i897_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i898_3_lut (.A(data_buffer_reg[905]), .B(\data_buffer[897] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[897])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i898_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i899_3_lut (.A(data_buffer_reg[906]), .B(\data_buffer[898] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[898])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i899_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i900_3_lut (.A(data_buffer_reg[907]), .B(\data_buffer[899] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[899])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i900_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i901_3_lut (.A(data_buffer_reg[908]), .B(\data_buffer[900] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[900])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i901_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i905_3_lut (.A(data_buffer_reg[912]), .B(\data_buffer[904] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[904])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i905_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i906_3_lut (.A(data_buffer_reg[913]), .B(\data_buffer[905] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[905])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i906_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i907_3_lut (.A(data_buffer_reg[914]), .B(\data_buffer[906] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[906])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i907_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i908_3_lut (.A(data_buffer_reg[915]), .B(\data_buffer[907] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[907])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i908_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i909_3_lut (.A(data_buffer_reg[916]), .B(\data_buffer[908] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[908])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i909_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i913_3_lut (.A(data_buffer_reg[920]), .B(\data_buffer[912] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[912])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i913_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i914_3_lut (.A(data_buffer_reg[921]), .B(\data_buffer[913] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[913])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i914_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i915_3_lut (.A(data_buffer_reg[922]), .B(\data_buffer[914] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[914])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i915_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i916_3_lut (.A(data_buffer_reg[923]), .B(\data_buffer[915] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[915])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i916_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i917_3_lut (.A(data_buffer_reg[924]), .B(\data_buffer[916] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[916])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i917_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i921_3_lut (.A(data_buffer_reg[928]), .B(\data_buffer[920] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[920])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i921_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i922_3_lut (.A(data_buffer_reg[929]), .B(\data_buffer[921] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[921])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i922_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i923_3_lut (.A(data_buffer_reg[930]), .B(\data_buffer[922] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[922])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i923_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_3_lut_4_lut_rep_488 (.A(data_length_reg[0]), .B(n15), 
         .C(n26793), .D(n25588), .Z(clk_c_enable_950)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i1_2_lut_3_lut_3_lut_4_lut_rep_488.init = 16'hfef0;
    LUT4 data_buffer_reg_959__I_0_i924_3_lut (.A(data_buffer_reg[931]), .B(\data_buffer[923] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[923])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i924_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i925_3_lut (.A(data_buffer_reg[932]), .B(\data_buffer[924] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[924])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i925_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i929_3_lut (.A(data_buffer_reg[936]), .B(\data_buffer[928] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[928])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i929_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i930_3_lut (.A(data_buffer_reg[937]), .B(\data_buffer[929] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[929])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i930_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i931_3_lut (.A(data_buffer_reg[938]), .B(\data_buffer[930] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[930])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i931_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i932_3_lut (.A(data_buffer_reg[939]), .B(\data_buffer[931] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[931])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i932_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i933_3_lut (.A(data_buffer_reg[940]), .B(\data_buffer[932] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[932])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i933_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i169_3_lut (.A(data_buffer_reg[176]), .B(\data_buffer[168] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[168])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i169_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i937_3_lut (.A(data_buffer_reg[944]), .B(\data_buffer[936] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[936])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i937_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i938_3_lut (.A(data_buffer_reg[945]), .B(\data_buffer[937] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[937])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i938_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i939_3_lut (.A(data_buffer_reg[946]), .B(\data_buffer[938] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[938])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i939_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i940_3_lut (.A(data_buffer_reg[947]), .B(\data_buffer[939] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[939])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i940_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i941_3_lut (.A(data_buffer_reg[948]), .B(\data_buffer[940] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[940])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i941_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i945_3_lut (.A(data_buffer_reg[952]), .B(\data_buffer[944] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[944])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i945_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i946_3_lut (.A(data_buffer_reg[953]), .B(\data_buffer[945] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[945])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i946_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i947_3_lut (.A(data_buffer_reg[954]), .B(\data_buffer[946] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[946])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i947_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i948_3_lut (.A(data_buffer_reg[955]), .B(\data_buffer[947] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[947])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i948_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i949_3_lut (.A(data_buffer_reg[956]), .B(\data_buffer[948] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[948])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i949_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_3_lut_4_lut_rep_489 (.A(data_length_reg[0]), .B(n15), 
         .C(n26793), .D(n25588), .Z(clk_c_enable_1000)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i1_2_lut_3_lut_3_lut_4_lut_rep_489.init = 16'hfef0;
    LUT4 i1_2_lut_3_lut_3_lut_4_lut_rep_493 (.A(data_length_reg[0]), .B(n15), 
         .C(n26793), .D(n25588), .Z(clk_c_enable_1200)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i1_2_lut_3_lut_3_lut_4_lut_rep_493.init = 16'hfef0;
    LUT4 data_buffer_reg_959__I_0_i170_3_lut (.A(data_buffer_reg[177]), .B(\data_buffer[169] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[169])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i170_3_lut.init = 16'hcaca;
    FD1P3AX data_buffer_reg_i1 (.D(data_buffer_reg_959__N_3020[1]), .SP(clk_c_enable_799), 
            .CK(clk_c), .Q(data_buffer_reg[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i1.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i2 (.D(data_buffer_reg_959__N_3020[2]), .SP(clk_c_enable_799), 
            .CK(clk_c), .Q(data_buffer_reg[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i2.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i3 (.D(data_buffer_reg_959__N_3020[3]), .SP(clk_c_enable_799), 
            .CK(clk_c), .Q(data_buffer_reg[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i3.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i4 (.D(data_buffer_reg_959__N_3020[4]), .SP(clk_c_enable_799), 
            .CK(clk_c), .Q(data_buffer_reg[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i4.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i8 (.D(data_buffer_reg_959__N_3020[8]), .SP(clk_c_enable_799), 
            .CK(clk_c), .Q(data_buffer_reg[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i8.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i9 (.D(data_buffer_reg_959__N_3020[9]), .SP(clk_c_enable_799), 
            .CK(clk_c), .Q(data_buffer_reg[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i9.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i10 (.D(data_buffer_reg_959__N_3020[10]), .SP(clk_c_enable_799), 
            .CK(clk_c), .Q(data_buffer_reg[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i10.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i11 (.D(data_buffer_reg_959__N_3020[11]), .SP(clk_c_enable_799), 
            .CK(clk_c), .Q(data_buffer_reg[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i11.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i12 (.D(data_buffer_reg_959__N_3020[12]), .SP(clk_c_enable_799), 
            .CK(clk_c), .Q(data_buffer_reg[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i12.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i16 (.D(data_buffer_reg_959__N_3020[16]), .SP(clk_c_enable_799), 
            .CK(clk_c), .Q(data_buffer_reg[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i16.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i17 (.D(data_buffer_reg_959__N_3020[17]), .SP(clk_c_enable_799), 
            .CK(clk_c), .Q(data_buffer_reg[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i17.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i18 (.D(data_buffer_reg_959__N_3020[18]), .SP(clk_c_enable_799), 
            .CK(clk_c), .Q(data_buffer_reg[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i18.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i19 (.D(data_buffer_reg_959__N_3020[19]), .SP(clk_c_enable_799), 
            .CK(clk_c), .Q(data_buffer_reg[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i19.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i20 (.D(data_buffer_reg_959__N_3020[20]), .SP(clk_c_enable_799), 
            .CK(clk_c), .Q(data_buffer_reg[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i20.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i24 (.D(data_buffer_reg_959__N_3020[24]), .SP(clk_c_enable_799), 
            .CK(clk_c), .Q(data_buffer_reg[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i24.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i25 (.D(data_buffer_reg_959__N_3020[25]), .SP(clk_c_enable_799), 
            .CK(clk_c), .Q(data_buffer_reg[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i25.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i26 (.D(data_buffer_reg_959__N_3020[26]), .SP(clk_c_enable_799), 
            .CK(clk_c), .Q(data_buffer_reg[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i26.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i27 (.D(data_buffer_reg_959__N_3020[27]), .SP(clk_c_enable_799), 
            .CK(clk_c), .Q(data_buffer_reg[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i27.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i28 (.D(data_buffer_reg_959__N_3020[28]), .SP(clk_c_enable_799), 
            .CK(clk_c), .Q(data_buffer_reg[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i28.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i32 (.D(data_buffer_reg_959__N_3020[32]), .SP(clk_c_enable_799), 
            .CK(clk_c), .Q(data_buffer_reg[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i32.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i33 (.D(data_buffer_reg_959__N_3020[33]), .SP(clk_c_enable_799), 
            .CK(clk_c), .Q(data_buffer_reg[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i33.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i34 (.D(data_buffer_reg_959__N_3020[34]), .SP(clk_c_enable_799), 
            .CK(clk_c), .Q(data_buffer_reg[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i34.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i35 (.D(data_buffer_reg_959__N_3020[35]), .SP(clk_c_enable_799), 
            .CK(clk_c), .Q(data_buffer_reg[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i35.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i36 (.D(data_buffer_reg_959__N_3020[36]), .SP(clk_c_enable_799), 
            .CK(clk_c), .Q(data_buffer_reg[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i36.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i40 (.D(data_buffer_reg_959__N_3020[40]), .SP(clk_c_enable_799), 
            .CK(clk_c), .Q(data_buffer_reg[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i40.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i41 (.D(data_buffer_reg_959__N_3020[41]), .SP(clk_c_enable_799), 
            .CK(clk_c), .Q(data_buffer_reg[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i41.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i42 (.D(data_buffer_reg_959__N_3020[42]), .SP(clk_c_enable_799), 
            .CK(clk_c), .Q(data_buffer_reg[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i42.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i43 (.D(data_buffer_reg_959__N_3020[43]), .SP(clk_c_enable_799), 
            .CK(clk_c), .Q(data_buffer_reg[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i43.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i44 (.D(data_buffer_reg_959__N_3020[44]), .SP(clk_c_enable_799), 
            .CK(clk_c), .Q(data_buffer_reg[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i44.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i48 (.D(data_buffer_reg_959__N_3020[48]), .SP(clk_c_enable_799), 
            .CK(clk_c), .Q(data_buffer_reg[48])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i48.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i49 (.D(data_buffer_reg_959__N_3020[49]), .SP(clk_c_enable_799), 
            .CK(clk_c), .Q(data_buffer_reg[49])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i49.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i50 (.D(data_buffer_reg_959__N_3020[50]), .SP(clk_c_enable_799), 
            .CK(clk_c), .Q(data_buffer_reg[50])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i50.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i51 (.D(data_buffer_reg_959__N_3020[51]), .SP(clk_c_enable_799), 
            .CK(clk_c), .Q(data_buffer_reg[51])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i51.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i52 (.D(data_buffer_reg_959__N_3020[52]), .SP(clk_c_enable_799), 
            .CK(clk_c), .Q(data_buffer_reg[52])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i52.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i56 (.D(data_buffer_reg_959__N_3020[56]), .SP(clk_c_enable_799), 
            .CK(clk_c), .Q(data_buffer_reg[56])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i56.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i57 (.D(data_buffer_reg_959__N_3020[57]), .SP(clk_c_enable_799), 
            .CK(clk_c), .Q(data_buffer_reg[57])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i57.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i58 (.D(data_buffer_reg_959__N_3020[58]), .SP(clk_c_enable_799), 
            .CK(clk_c), .Q(data_buffer_reg[58])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i58.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i59 (.D(data_buffer_reg_959__N_3020[59]), .SP(clk_c_enable_799), 
            .CK(clk_c), .Q(data_buffer_reg[59])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i59.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i60 (.D(data_buffer_reg_959__N_3020[60]), .SP(clk_c_enable_799), 
            .CK(clk_c), .Q(data_buffer_reg[60])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i60.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i64 (.D(data_buffer_reg_959__N_3020[64]), .SP(clk_c_enable_799), 
            .CK(clk_c), .Q(data_buffer_reg[64])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i64.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i65 (.D(data_buffer_reg_959__N_3020[65]), .SP(clk_c_enable_799), 
            .CK(clk_c), .Q(data_buffer_reg[65])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i65.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i66 (.D(data_buffer_reg_959__N_3020[66]), .SP(clk_c_enable_799), 
            .CK(clk_c), .Q(data_buffer_reg[66])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i66.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i67 (.D(data_buffer_reg_959__N_3020[67]), .SP(clk_c_enable_799), 
            .CK(clk_c), .Q(data_buffer_reg[67])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i67.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i68 (.D(data_buffer_reg_959__N_3020[68]), .SP(clk_c_enable_799), 
            .CK(clk_c), .Q(data_buffer_reg[68])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i68.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i72 (.D(data_buffer_reg_959__N_3020[72]), .SP(clk_c_enable_799), 
            .CK(clk_c), .Q(data_buffer_reg[72])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i72.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i73 (.D(data_buffer_reg_959__N_3020[73]), .SP(clk_c_enable_799), 
            .CK(clk_c), .Q(data_buffer_reg[73])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i73.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i74 (.D(data_buffer_reg_959__N_3020[74]), .SP(clk_c_enable_799), 
            .CK(clk_c), .Q(data_buffer_reg[74])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i74.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i75 (.D(data_buffer_reg_959__N_3020[75]), .SP(clk_c_enable_799), 
            .CK(clk_c), .Q(data_buffer_reg[75])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i75.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i76 (.D(data_buffer_reg_959__N_3020[76]), .SP(clk_c_enable_799), 
            .CK(clk_c), .Q(data_buffer_reg[76])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i76.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i80 (.D(data_buffer_reg_959__N_3020[80]), .SP(clk_c_enable_849), 
            .CK(clk_c), .Q(data_buffer_reg[80])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i80.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i81 (.D(data_buffer_reg_959__N_3020[81]), .SP(clk_c_enable_849), 
            .CK(clk_c), .Q(data_buffer_reg[81])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i81.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i82 (.D(data_buffer_reg_959__N_3020[82]), .SP(clk_c_enable_849), 
            .CK(clk_c), .Q(data_buffer_reg[82])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i82.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i83 (.D(data_buffer_reg_959__N_3020[83]), .SP(clk_c_enable_849), 
            .CK(clk_c), .Q(data_buffer_reg[83])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i83.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i84 (.D(data_buffer_reg_959__N_3020[84]), .SP(clk_c_enable_849), 
            .CK(clk_c), .Q(data_buffer_reg[84])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i84.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i88 (.D(data_buffer_reg_959__N_3020[88]), .SP(clk_c_enable_849), 
            .CK(clk_c), .Q(data_buffer_reg[88])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i88.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i89 (.D(data_buffer_reg_959__N_3020[89]), .SP(clk_c_enable_849), 
            .CK(clk_c), .Q(data_buffer_reg[89])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i89.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i90 (.D(data_buffer_reg_959__N_3020[90]), .SP(clk_c_enable_849), 
            .CK(clk_c), .Q(data_buffer_reg[90])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i90.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i91 (.D(data_buffer_reg_959__N_3020[91]), .SP(clk_c_enable_849), 
            .CK(clk_c), .Q(data_buffer_reg[91])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i91.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i92 (.D(data_buffer_reg_959__N_3020[92]), .SP(clk_c_enable_849), 
            .CK(clk_c), .Q(data_buffer_reg[92])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i92.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i96 (.D(data_buffer_reg_959__N_3020[96]), .SP(clk_c_enable_849), 
            .CK(clk_c), .Q(data_buffer_reg[96])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i96.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i97 (.D(data_buffer_reg_959__N_3020[97]), .SP(clk_c_enable_849), 
            .CK(clk_c), .Q(data_buffer_reg[97])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i97.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i98 (.D(data_buffer_reg_959__N_3020[98]), .SP(clk_c_enable_849), 
            .CK(clk_c), .Q(data_buffer_reg[98])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i98.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i99 (.D(data_buffer_reg_959__N_3020[99]), .SP(clk_c_enable_849), 
            .CK(clk_c), .Q(data_buffer_reg[99])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i99.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i100 (.D(data_buffer_reg_959__N_3020[100]), .SP(clk_c_enable_849), 
            .CK(clk_c), .Q(data_buffer_reg[100])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i100.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i104 (.D(data_buffer_reg_959__N_3020[104]), .SP(clk_c_enable_849), 
            .CK(clk_c), .Q(data_buffer_reg[104])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i104.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i105 (.D(data_buffer_reg_959__N_3020[105]), .SP(clk_c_enable_849), 
            .CK(clk_c), .Q(data_buffer_reg[105])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i105.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i106 (.D(data_buffer_reg_959__N_3020[106]), .SP(clk_c_enable_849), 
            .CK(clk_c), .Q(data_buffer_reg[106])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i106.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i107 (.D(data_buffer_reg_959__N_3020[107]), .SP(clk_c_enable_849), 
            .CK(clk_c), .Q(data_buffer_reg[107])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i107.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i108 (.D(data_buffer_reg_959__N_3020[108]), .SP(clk_c_enable_849), 
            .CK(clk_c), .Q(data_buffer_reg[108])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i108.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i112 (.D(data_buffer_reg_959__N_3020[112]), .SP(clk_c_enable_849), 
            .CK(clk_c), .Q(data_buffer_reg[112])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i112.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i113 (.D(data_buffer_reg_959__N_3020[113]), .SP(clk_c_enable_849), 
            .CK(clk_c), .Q(data_buffer_reg[113])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i113.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i114 (.D(data_buffer_reg_959__N_3020[114]), .SP(clk_c_enable_849), 
            .CK(clk_c), .Q(data_buffer_reg[114])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i114.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i115 (.D(data_buffer_reg_959__N_3020[115]), .SP(clk_c_enable_849), 
            .CK(clk_c), .Q(data_buffer_reg[115])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i115.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i116 (.D(data_buffer_reg_959__N_3020[116]), .SP(clk_c_enable_849), 
            .CK(clk_c), .Q(data_buffer_reg[116])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i116.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i120 (.D(data_buffer_reg_959__N_3020[120]), .SP(clk_c_enable_849), 
            .CK(clk_c), .Q(data_buffer_reg[120])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i120.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i121 (.D(data_buffer_reg_959__N_3020[121]), .SP(clk_c_enable_849), 
            .CK(clk_c), .Q(data_buffer_reg[121])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i121.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i122 (.D(data_buffer_reg_959__N_3020[122]), .SP(clk_c_enable_849), 
            .CK(clk_c), .Q(data_buffer_reg[122])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i122.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i123 (.D(data_buffer_reg_959__N_3020[123]), .SP(clk_c_enable_849), 
            .CK(clk_c), .Q(data_buffer_reg[123])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i123.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i124 (.D(data_buffer_reg_959__N_3020[124]), .SP(clk_c_enable_849), 
            .CK(clk_c), .Q(data_buffer_reg[124])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i124.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i128 (.D(data_buffer_reg_959__N_3020[128]), .SP(clk_c_enable_849), 
            .CK(clk_c), .Q(data_buffer_reg[128])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i128.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i129 (.D(data_buffer_reg_959__N_3020[129]), .SP(clk_c_enable_849), 
            .CK(clk_c), .Q(data_buffer_reg[129])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i129.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i130 (.D(data_buffer_reg_959__N_3020[130]), .SP(clk_c_enable_849), 
            .CK(clk_c), .Q(data_buffer_reg[130])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i130.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i131 (.D(data_buffer_reg_959__N_3020[131]), .SP(clk_c_enable_849), 
            .CK(clk_c), .Q(data_buffer_reg[131])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i131.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i132 (.D(data_buffer_reg_959__N_3020[132]), .SP(clk_c_enable_849), 
            .CK(clk_c), .Q(data_buffer_reg[132])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i132.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i136 (.D(data_buffer_reg_959__N_3020[136]), .SP(clk_c_enable_849), 
            .CK(clk_c), .Q(data_buffer_reg[136])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i136.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i137 (.D(data_buffer_reg_959__N_3020[137]), .SP(clk_c_enable_849), 
            .CK(clk_c), .Q(data_buffer_reg[137])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i137.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i138 (.D(data_buffer_reg_959__N_3020[138]), .SP(clk_c_enable_849), 
            .CK(clk_c), .Q(data_buffer_reg[138])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i138.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i139 (.D(data_buffer_reg_959__N_3020[139]), .SP(clk_c_enable_849), 
            .CK(clk_c), .Q(data_buffer_reg[139])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i139.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i140 (.D(data_buffer_reg_959__N_3020[140]), .SP(clk_c_enable_849), 
            .CK(clk_c), .Q(data_buffer_reg[140])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i140.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i144 (.D(data_buffer_reg_959__N_3020[144]), .SP(clk_c_enable_849), 
            .CK(clk_c), .Q(data_buffer_reg[144])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i144.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i145 (.D(data_buffer_reg_959__N_3020[145]), .SP(clk_c_enable_849), 
            .CK(clk_c), .Q(data_buffer_reg[145])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i145.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i146 (.D(data_buffer_reg_959__N_3020[146]), .SP(clk_c_enable_849), 
            .CK(clk_c), .Q(data_buffer_reg[146])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i146.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i147 (.D(data_buffer_reg_959__N_3020[147]), .SP(clk_c_enable_849), 
            .CK(clk_c), .Q(data_buffer_reg[147])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i147.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i148 (.D(data_buffer_reg_959__N_3020[148]), .SP(clk_c_enable_849), 
            .CK(clk_c), .Q(data_buffer_reg[148])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i148.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i152 (.D(data_buffer_reg_959__N_3020[152]), .SP(clk_c_enable_849), 
            .CK(clk_c), .Q(data_buffer_reg[152])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i152.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i153 (.D(data_buffer_reg_959__N_3020[153]), .SP(clk_c_enable_849), 
            .CK(clk_c), .Q(data_buffer_reg[153])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i153.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i154 (.D(data_buffer_reg_959__N_3020[154]), .SP(clk_c_enable_849), 
            .CK(clk_c), .Q(data_buffer_reg[154])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i154.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i155 (.D(data_buffer_reg_959__N_3020[155]), .SP(clk_c_enable_849), 
            .CK(clk_c), .Q(data_buffer_reg[155])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i155.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i156 (.D(data_buffer_reg_959__N_3020[156]), .SP(clk_c_enable_849), 
            .CK(clk_c), .Q(data_buffer_reg[156])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i156.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i160 (.D(data_buffer_reg_959__N_3020[160]), .SP(clk_c_enable_899), 
            .CK(clk_c), .Q(data_buffer_reg[160])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i160.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i161 (.D(data_buffer_reg_959__N_3020[161]), .SP(clk_c_enable_899), 
            .CK(clk_c), .Q(data_buffer_reg[161])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i161.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i162 (.D(data_buffer_reg_959__N_3020[162]), .SP(clk_c_enable_899), 
            .CK(clk_c), .Q(data_buffer_reg[162])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i162.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i163 (.D(data_buffer_reg_959__N_3020[163]), .SP(clk_c_enable_899), 
            .CK(clk_c), .Q(data_buffer_reg[163])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i163.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i164 (.D(data_buffer_reg_959__N_3020[164]), .SP(clk_c_enable_899), 
            .CK(clk_c), .Q(data_buffer_reg[164])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i164.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i168 (.D(data_buffer_reg_959__N_3020[168]), .SP(clk_c_enable_899), 
            .CK(clk_c), .Q(data_buffer_reg[168])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i168.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i169 (.D(data_buffer_reg_959__N_3020[169]), .SP(clk_c_enable_899), 
            .CK(clk_c), .Q(data_buffer_reg[169])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i169.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i170 (.D(data_buffer_reg_959__N_3020[170]), .SP(clk_c_enable_899), 
            .CK(clk_c), .Q(data_buffer_reg[170])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i170.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i171 (.D(data_buffer_reg_959__N_3020[171]), .SP(clk_c_enable_899), 
            .CK(clk_c), .Q(data_buffer_reg[171])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i171.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i172 (.D(data_buffer_reg_959__N_3020[172]), .SP(clk_c_enable_899), 
            .CK(clk_c), .Q(data_buffer_reg[172])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i172.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i176 (.D(data_buffer_reg_959__N_3020[176]), .SP(clk_c_enable_899), 
            .CK(clk_c), .Q(data_buffer_reg[176])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i176.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i177 (.D(data_buffer_reg_959__N_3020[177]), .SP(clk_c_enable_899), 
            .CK(clk_c), .Q(data_buffer_reg[177])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i177.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i178 (.D(data_buffer_reg_959__N_3020[178]), .SP(clk_c_enable_899), 
            .CK(clk_c), .Q(data_buffer_reg[178])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i178.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i179 (.D(data_buffer_reg_959__N_3020[179]), .SP(clk_c_enable_899), 
            .CK(clk_c), .Q(data_buffer_reg[179])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i179.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i180 (.D(data_buffer_reg_959__N_3020[180]), .SP(clk_c_enable_899), 
            .CK(clk_c), .Q(data_buffer_reg[180])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i180.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i184 (.D(data_buffer_reg_959__N_3020[184]), .SP(clk_c_enable_899), 
            .CK(clk_c), .Q(data_buffer_reg[184])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i184.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i185 (.D(data_buffer_reg_959__N_3020[185]), .SP(clk_c_enable_899), 
            .CK(clk_c), .Q(data_buffer_reg[185])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i185.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i186 (.D(data_buffer_reg_959__N_3020[186]), .SP(clk_c_enable_899), 
            .CK(clk_c), .Q(data_buffer_reg[186])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i186.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i187 (.D(data_buffer_reg_959__N_3020[187]), .SP(clk_c_enable_899), 
            .CK(clk_c), .Q(data_buffer_reg[187])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i187.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i188 (.D(data_buffer_reg_959__N_3020[188]), .SP(clk_c_enable_899), 
            .CK(clk_c), .Q(data_buffer_reg[188])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i188.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i192 (.D(data_buffer_reg_959__N_3020[192]), .SP(clk_c_enable_899), 
            .CK(clk_c), .Q(data_buffer_reg[192])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i192.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i193 (.D(data_buffer_reg_959__N_3020[193]), .SP(clk_c_enable_899), 
            .CK(clk_c), .Q(data_buffer_reg[193])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i193.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i194 (.D(data_buffer_reg_959__N_3020[194]), .SP(clk_c_enable_899), 
            .CK(clk_c), .Q(data_buffer_reg[194])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i194.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i195 (.D(data_buffer_reg_959__N_3020[195]), .SP(clk_c_enable_899), 
            .CK(clk_c), .Q(data_buffer_reg[195])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i195.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i196 (.D(data_buffer_reg_959__N_3020[196]), .SP(clk_c_enable_899), 
            .CK(clk_c), .Q(data_buffer_reg[196])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i196.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i200 (.D(data_buffer_reg_959__N_3020[200]), .SP(clk_c_enable_899), 
            .CK(clk_c), .Q(data_buffer_reg[200])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i200.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i201 (.D(data_buffer_reg_959__N_3020[201]), .SP(clk_c_enable_899), 
            .CK(clk_c), .Q(data_buffer_reg[201])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i201.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i202 (.D(data_buffer_reg_959__N_3020[202]), .SP(clk_c_enable_899), 
            .CK(clk_c), .Q(data_buffer_reg[202])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i202.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i203 (.D(data_buffer_reg_959__N_3020[203]), .SP(clk_c_enable_899), 
            .CK(clk_c), .Q(data_buffer_reg[203])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i203.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i204 (.D(data_buffer_reg_959__N_3020[204]), .SP(clk_c_enable_899), 
            .CK(clk_c), .Q(data_buffer_reg[204])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i204.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i208 (.D(data_buffer_reg_959__N_3020[208]), .SP(clk_c_enable_899), 
            .CK(clk_c), .Q(data_buffer_reg[208])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i208.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i209 (.D(data_buffer_reg_959__N_3020[209]), .SP(clk_c_enable_899), 
            .CK(clk_c), .Q(data_buffer_reg[209])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i209.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i210 (.D(data_buffer_reg_959__N_3020[210]), .SP(clk_c_enable_899), 
            .CK(clk_c), .Q(data_buffer_reg[210])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i210.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i211 (.D(data_buffer_reg_959__N_3020[211]), .SP(clk_c_enable_899), 
            .CK(clk_c), .Q(data_buffer_reg[211])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i211.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i212 (.D(data_buffer_reg_959__N_3020[212]), .SP(clk_c_enable_899), 
            .CK(clk_c), .Q(data_buffer_reg[212])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i212.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i216 (.D(data_buffer_reg_959__N_3020[216]), .SP(clk_c_enable_899), 
            .CK(clk_c), .Q(data_buffer_reg[216])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i216.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i217 (.D(data_buffer_reg_959__N_3020[217]), .SP(clk_c_enable_899), 
            .CK(clk_c), .Q(data_buffer_reg[217])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i217.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i218 (.D(data_buffer_reg_959__N_3020[218]), .SP(clk_c_enable_899), 
            .CK(clk_c), .Q(data_buffer_reg[218])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i218.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i219 (.D(data_buffer_reg_959__N_3020[219]), .SP(clk_c_enable_899), 
            .CK(clk_c), .Q(data_buffer_reg[219])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i219.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i220 (.D(data_buffer_reg_959__N_3020[220]), .SP(clk_c_enable_899), 
            .CK(clk_c), .Q(data_buffer_reg[220])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i220.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i224 (.D(data_buffer_reg_959__N_3020[224]), .SP(clk_c_enable_899), 
            .CK(clk_c), .Q(data_buffer_reg[224])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i224.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i225 (.D(data_buffer_reg_959__N_3020[225]), .SP(clk_c_enable_899), 
            .CK(clk_c), .Q(data_buffer_reg[225])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i225.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i226 (.D(data_buffer_reg_959__N_3020[226]), .SP(clk_c_enable_899), 
            .CK(clk_c), .Q(data_buffer_reg[226])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i226.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i227 (.D(data_buffer_reg_959__N_3020[227]), .SP(clk_c_enable_899), 
            .CK(clk_c), .Q(data_buffer_reg[227])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i227.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i228 (.D(data_buffer_reg_959__N_3020[228]), .SP(clk_c_enable_899), 
            .CK(clk_c), .Q(data_buffer_reg[228])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i228.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i232 (.D(data_buffer_reg_959__N_3020[232]), .SP(clk_c_enable_899), 
            .CK(clk_c), .Q(data_buffer_reg[232])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i232.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i233 (.D(data_buffer_reg_959__N_3020[233]), .SP(clk_c_enable_899), 
            .CK(clk_c), .Q(data_buffer_reg[233])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i233.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i234 (.D(data_buffer_reg_959__N_3020[234]), .SP(clk_c_enable_899), 
            .CK(clk_c), .Q(data_buffer_reg[234])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i234.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i235 (.D(data_buffer_reg_959__N_3020[235]), .SP(clk_c_enable_899), 
            .CK(clk_c), .Q(data_buffer_reg[235])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i235.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i236 (.D(data_buffer_reg_959__N_3020[236]), .SP(clk_c_enable_899), 
            .CK(clk_c), .Q(data_buffer_reg[236])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i236.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i240 (.D(data_buffer_reg_959__N_3020[240]), .SP(clk_c_enable_950), 
            .CK(clk_c), .Q(data_buffer_reg[240])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i240.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i241 (.D(data_buffer_reg_959__N_3020[241]), .SP(clk_c_enable_950), 
            .CK(clk_c), .Q(data_buffer_reg[241])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i241.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i242 (.D(data_buffer_reg_959__N_3020[242]), .SP(clk_c_enable_950), 
            .CK(clk_c), .Q(data_buffer_reg[242])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i242.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i243 (.D(data_buffer_reg_959__N_3020[243]), .SP(clk_c_enable_950), 
            .CK(clk_c), .Q(data_buffer_reg[243])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i243.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i244 (.D(data_buffer_reg_959__N_3020[244]), .SP(clk_c_enable_950), 
            .CK(clk_c), .Q(data_buffer_reg[244])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i244.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i248 (.D(data_buffer_reg_959__N_3020[248]), .SP(clk_c_enable_950), 
            .CK(clk_c), .Q(data_buffer_reg[248])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i248.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i249 (.D(data_buffer_reg_959__N_3020[249]), .SP(clk_c_enable_950), 
            .CK(clk_c), .Q(data_buffer_reg[249])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i249.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i250 (.D(data_buffer_reg_959__N_3020[250]), .SP(clk_c_enable_950), 
            .CK(clk_c), .Q(data_buffer_reg[250])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i250.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i251 (.D(data_buffer_reg_959__N_3020[251]), .SP(clk_c_enable_950), 
            .CK(clk_c), .Q(data_buffer_reg[251])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i251.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i252 (.D(data_buffer_reg_959__N_3020[252]), .SP(clk_c_enable_950), 
            .CK(clk_c), .Q(data_buffer_reg[252])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i252.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i256 (.D(data_buffer_reg_959__N_3020[256]), .SP(clk_c_enable_950), 
            .CK(clk_c), .Q(data_buffer_reg[256])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i256.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i257 (.D(data_buffer_reg_959__N_3020[257]), .SP(clk_c_enable_950), 
            .CK(clk_c), .Q(data_buffer_reg[257])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i257.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i258 (.D(data_buffer_reg_959__N_3020[258]), .SP(clk_c_enable_950), 
            .CK(clk_c), .Q(data_buffer_reg[258])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i258.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i259 (.D(data_buffer_reg_959__N_3020[259]), .SP(clk_c_enable_950), 
            .CK(clk_c), .Q(data_buffer_reg[259])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i259.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i260 (.D(data_buffer_reg_959__N_3020[260]), .SP(clk_c_enable_950), 
            .CK(clk_c), .Q(data_buffer_reg[260])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i260.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i264 (.D(data_buffer_reg_959__N_3020[264]), .SP(clk_c_enable_950), 
            .CK(clk_c), .Q(data_buffer_reg[264])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i264.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i265 (.D(data_buffer_reg_959__N_3020[265]), .SP(clk_c_enable_950), 
            .CK(clk_c), .Q(data_buffer_reg[265])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i265.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i266 (.D(data_buffer_reg_959__N_3020[266]), .SP(clk_c_enable_950), 
            .CK(clk_c), .Q(data_buffer_reg[266])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i266.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i267 (.D(data_buffer_reg_959__N_3020[267]), .SP(clk_c_enable_950), 
            .CK(clk_c), .Q(data_buffer_reg[267])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i267.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i268 (.D(data_buffer_reg_959__N_3020[268]), .SP(clk_c_enable_950), 
            .CK(clk_c), .Q(data_buffer_reg[268])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i268.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i272 (.D(data_buffer_reg_959__N_3020[272]), .SP(clk_c_enable_950), 
            .CK(clk_c), .Q(data_buffer_reg[272])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i272.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i273 (.D(data_buffer_reg_959__N_3020[273]), .SP(clk_c_enable_950), 
            .CK(clk_c), .Q(data_buffer_reg[273])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i273.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i274 (.D(data_buffer_reg_959__N_3020[274]), .SP(clk_c_enable_950), 
            .CK(clk_c), .Q(data_buffer_reg[274])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i274.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i275 (.D(data_buffer_reg_959__N_3020[275]), .SP(clk_c_enable_950), 
            .CK(clk_c), .Q(data_buffer_reg[275])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i275.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i276 (.D(data_buffer_reg_959__N_3020[276]), .SP(clk_c_enable_950), 
            .CK(clk_c), .Q(data_buffer_reg[276])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i276.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i280 (.D(data_buffer_reg_959__N_3020[280]), .SP(clk_c_enable_950), 
            .CK(clk_c), .Q(data_buffer_reg[280])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i280.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i281 (.D(data_buffer_reg_959__N_3020[281]), .SP(clk_c_enable_950), 
            .CK(clk_c), .Q(data_buffer_reg[281])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i281.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i282 (.D(data_buffer_reg_959__N_3020[282]), .SP(clk_c_enable_950), 
            .CK(clk_c), .Q(data_buffer_reg[282])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i282.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i283 (.D(data_buffer_reg_959__N_3020[283]), .SP(clk_c_enable_950), 
            .CK(clk_c), .Q(data_buffer_reg[283])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i283.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i284 (.D(data_buffer_reg_959__N_3020[284]), .SP(clk_c_enable_950), 
            .CK(clk_c), .Q(data_buffer_reg[284])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i284.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i288 (.D(data_buffer_reg_959__N_3020[288]), .SP(clk_c_enable_950), 
            .CK(clk_c), .Q(data_buffer_reg[288])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i288.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i289 (.D(data_buffer_reg_959__N_3020[289]), .SP(clk_c_enable_950), 
            .CK(clk_c), .Q(data_buffer_reg[289])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i289.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i290 (.D(data_buffer_reg_959__N_3020[290]), .SP(clk_c_enable_950), 
            .CK(clk_c), .Q(data_buffer_reg[290])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i290.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i291 (.D(data_buffer_reg_959__N_3020[291]), .SP(clk_c_enable_950), 
            .CK(clk_c), .Q(data_buffer_reg[291])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i291.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i292 (.D(data_buffer_reg_959__N_3020[292]), .SP(clk_c_enable_950), 
            .CK(clk_c), .Q(data_buffer_reg[292])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i292.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i296 (.D(data_buffer_reg_959__N_3020[296]), .SP(clk_c_enable_950), 
            .CK(clk_c), .Q(data_buffer_reg[296])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i296.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i297 (.D(data_buffer_reg_959__N_3020[297]), .SP(clk_c_enable_950), 
            .CK(clk_c), .Q(data_buffer_reg[297])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i297.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i298 (.D(data_buffer_reg_959__N_3020[298]), .SP(clk_c_enable_950), 
            .CK(clk_c), .Q(data_buffer_reg[298])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i298.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i299 (.D(data_buffer_reg_959__N_3020[299]), .SP(clk_c_enable_950), 
            .CK(clk_c), .Q(data_buffer_reg[299])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i299.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i300 (.D(data_buffer_reg_959__N_3020[300]), .SP(clk_c_enable_950), 
            .CK(clk_c), .Q(data_buffer_reg[300])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i300.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i304 (.D(data_buffer_reg_959__N_3020[304]), .SP(clk_c_enable_950), 
            .CK(clk_c), .Q(data_buffer_reg[304])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i304.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i305 (.D(data_buffer_reg_959__N_3020[305]), .SP(clk_c_enable_950), 
            .CK(clk_c), .Q(data_buffer_reg[305])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i305.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i306 (.D(data_buffer_reg_959__N_3020[306]), .SP(clk_c_enable_950), 
            .CK(clk_c), .Q(data_buffer_reg[306])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i306.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i307 (.D(data_buffer_reg_959__N_3020[307]), .SP(clk_c_enable_950), 
            .CK(clk_c), .Q(data_buffer_reg[307])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i307.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i308 (.D(data_buffer_reg_959__N_3020[308]), .SP(clk_c_enable_950), 
            .CK(clk_c), .Q(data_buffer_reg[308])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i308.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i312 (.D(data_buffer_reg_959__N_3020[312]), .SP(clk_c_enable_950), 
            .CK(clk_c), .Q(data_buffer_reg[312])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i312.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i313 (.D(data_buffer_reg_959__N_3020[313]), .SP(clk_c_enable_950), 
            .CK(clk_c), .Q(data_buffer_reg[313])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i313.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i314 (.D(data_buffer_reg_959__N_3020[314]), .SP(clk_c_enable_950), 
            .CK(clk_c), .Q(data_buffer_reg[314])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i314.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i315 (.D(data_buffer_reg_959__N_3020[315]), .SP(clk_c_enable_950), 
            .CK(clk_c), .Q(data_buffer_reg[315])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i315.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i316 (.D(data_buffer_reg_959__N_3020[316]), .SP(clk_c_enable_950), 
            .CK(clk_c), .Q(data_buffer_reg[316])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i316.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i320 (.D(data_buffer_reg_959__N_3020[320]), .SP(clk_c_enable_1000), 
            .CK(clk_c), .Q(data_buffer_reg[320])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i320.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i321 (.D(data_buffer_reg_959__N_3020[321]), .SP(clk_c_enable_1000), 
            .CK(clk_c), .Q(data_buffer_reg[321])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i321.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i322 (.D(data_buffer_reg_959__N_3020[322]), .SP(clk_c_enable_1000), 
            .CK(clk_c), .Q(data_buffer_reg[322])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i322.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i323 (.D(data_buffer_reg_959__N_3020[323]), .SP(clk_c_enable_1000), 
            .CK(clk_c), .Q(data_buffer_reg[323])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i323.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i324 (.D(data_buffer_reg_959__N_3020[324]), .SP(clk_c_enable_1000), 
            .CK(clk_c), .Q(data_buffer_reg[324])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i324.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i328 (.D(data_buffer_reg_959__N_3020[328]), .SP(clk_c_enable_1000), 
            .CK(clk_c), .Q(data_buffer_reg[328])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i328.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i329 (.D(data_buffer_reg_959__N_3020[329]), .SP(clk_c_enable_1000), 
            .CK(clk_c), .Q(data_buffer_reg[329])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i329.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i330 (.D(data_buffer_reg_959__N_3020[330]), .SP(clk_c_enable_1000), 
            .CK(clk_c), .Q(data_buffer_reg[330])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i330.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i331 (.D(data_buffer_reg_959__N_3020[331]), .SP(clk_c_enable_1000), 
            .CK(clk_c), .Q(data_buffer_reg[331])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i331.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i332 (.D(data_buffer_reg_959__N_3020[332]), .SP(clk_c_enable_1000), 
            .CK(clk_c), .Q(data_buffer_reg[332])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i332.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i336 (.D(data_buffer_reg_959__N_3020[336]), .SP(clk_c_enable_1000), 
            .CK(clk_c), .Q(data_buffer_reg[336])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i336.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i337 (.D(data_buffer_reg_959__N_3020[337]), .SP(clk_c_enable_1000), 
            .CK(clk_c), .Q(data_buffer_reg[337])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i337.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i338 (.D(data_buffer_reg_959__N_3020[338]), .SP(clk_c_enable_1000), 
            .CK(clk_c), .Q(data_buffer_reg[338])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i338.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i339 (.D(data_buffer_reg_959__N_3020[339]), .SP(clk_c_enable_1000), 
            .CK(clk_c), .Q(data_buffer_reg[339])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i339.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i340 (.D(data_buffer_reg_959__N_3020[340]), .SP(clk_c_enable_1000), 
            .CK(clk_c), .Q(data_buffer_reg[340])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i340.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i344 (.D(data_buffer_reg_959__N_3020[344]), .SP(clk_c_enable_1000), 
            .CK(clk_c), .Q(data_buffer_reg[344])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i344.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i345 (.D(data_buffer_reg_959__N_3020[345]), .SP(clk_c_enable_1000), 
            .CK(clk_c), .Q(data_buffer_reg[345])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i345.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i346 (.D(data_buffer_reg_959__N_3020[346]), .SP(clk_c_enable_1000), 
            .CK(clk_c), .Q(data_buffer_reg[346])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i346.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i347 (.D(data_buffer_reg_959__N_3020[347]), .SP(clk_c_enable_1000), 
            .CK(clk_c), .Q(data_buffer_reg[347])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i347.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i348 (.D(data_buffer_reg_959__N_3020[348]), .SP(clk_c_enable_1000), 
            .CK(clk_c), .Q(data_buffer_reg[348])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i348.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i352 (.D(data_buffer_reg_959__N_3020[352]), .SP(clk_c_enable_1000), 
            .CK(clk_c), .Q(data_buffer_reg[352])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i352.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i353 (.D(data_buffer_reg_959__N_3020[353]), .SP(clk_c_enable_1000), 
            .CK(clk_c), .Q(data_buffer_reg[353])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i353.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i354 (.D(data_buffer_reg_959__N_3020[354]), .SP(clk_c_enable_1000), 
            .CK(clk_c), .Q(data_buffer_reg[354])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i354.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i355 (.D(data_buffer_reg_959__N_3020[355]), .SP(clk_c_enable_1000), 
            .CK(clk_c), .Q(data_buffer_reg[355])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i355.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i356 (.D(data_buffer_reg_959__N_3020[356]), .SP(clk_c_enable_1000), 
            .CK(clk_c), .Q(data_buffer_reg[356])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i356.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i360 (.D(data_buffer_reg_959__N_3020[360]), .SP(clk_c_enable_1000), 
            .CK(clk_c), .Q(data_buffer_reg[360])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i360.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i361 (.D(data_buffer_reg_959__N_3020[361]), .SP(clk_c_enable_1000), 
            .CK(clk_c), .Q(data_buffer_reg[361])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i361.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i362 (.D(data_buffer_reg_959__N_3020[362]), .SP(clk_c_enable_1000), 
            .CK(clk_c), .Q(data_buffer_reg[362])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i362.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i363 (.D(data_buffer_reg_959__N_3020[363]), .SP(clk_c_enable_1000), 
            .CK(clk_c), .Q(data_buffer_reg[363])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i363.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i364 (.D(data_buffer_reg_959__N_3020[364]), .SP(clk_c_enable_1000), 
            .CK(clk_c), .Q(data_buffer_reg[364])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i364.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i368 (.D(data_buffer_reg_959__N_3020[368]), .SP(clk_c_enable_1000), 
            .CK(clk_c), .Q(data_buffer_reg[368])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i368.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i369 (.D(data_buffer_reg_959__N_3020[369]), .SP(clk_c_enable_1000), 
            .CK(clk_c), .Q(data_buffer_reg[369])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i369.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i370 (.D(data_buffer_reg_959__N_3020[370]), .SP(clk_c_enable_1000), 
            .CK(clk_c), .Q(data_buffer_reg[370])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i370.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i371 (.D(data_buffer_reg_959__N_3020[371]), .SP(clk_c_enable_1000), 
            .CK(clk_c), .Q(data_buffer_reg[371])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i371.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i372 (.D(data_buffer_reg_959__N_3020[372]), .SP(clk_c_enable_1000), 
            .CK(clk_c), .Q(data_buffer_reg[372])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i372.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i376 (.D(data_buffer_reg_959__N_3020[376]), .SP(clk_c_enable_1000), 
            .CK(clk_c), .Q(data_buffer_reg[376])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i376.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i377 (.D(data_buffer_reg_959__N_3020[377]), .SP(clk_c_enable_1000), 
            .CK(clk_c), .Q(data_buffer_reg[377])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i377.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i378 (.D(data_buffer_reg_959__N_3020[378]), .SP(clk_c_enable_1000), 
            .CK(clk_c), .Q(data_buffer_reg[378])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i378.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i379 (.D(data_buffer_reg_959__N_3020[379]), .SP(clk_c_enable_1000), 
            .CK(clk_c), .Q(data_buffer_reg[379])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i379.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i380 (.D(data_buffer_reg_959__N_3020[380]), .SP(clk_c_enable_1000), 
            .CK(clk_c), .Q(data_buffer_reg[380])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i380.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i384 (.D(data_buffer_reg_959__N_3020[384]), .SP(clk_c_enable_1000), 
            .CK(clk_c), .Q(data_buffer_reg[384])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i384.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i385 (.D(data_buffer_reg_959__N_3020[385]), .SP(clk_c_enable_1000), 
            .CK(clk_c), .Q(data_buffer_reg[385])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i385.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i386 (.D(data_buffer_reg_959__N_3020[386]), .SP(clk_c_enable_1000), 
            .CK(clk_c), .Q(data_buffer_reg[386])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i386.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i387 (.D(data_buffer_reg_959__N_3020[387]), .SP(clk_c_enable_1000), 
            .CK(clk_c), .Q(data_buffer_reg[387])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i387.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i388 (.D(data_buffer_reg_959__N_3020[388]), .SP(clk_c_enable_1000), 
            .CK(clk_c), .Q(data_buffer_reg[388])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i388.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i392 (.D(data_buffer_reg_959__N_3020[392]), .SP(clk_c_enable_1000), 
            .CK(clk_c), .Q(data_buffer_reg[392])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i392.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i393 (.D(data_buffer_reg_959__N_3020[393]), .SP(clk_c_enable_1000), 
            .CK(clk_c), .Q(data_buffer_reg[393])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i393.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i394 (.D(data_buffer_reg_959__N_3020[394]), .SP(clk_c_enable_1000), 
            .CK(clk_c), .Q(data_buffer_reg[394])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i394.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i395 (.D(data_buffer_reg_959__N_3020[395]), .SP(clk_c_enable_1000), 
            .CK(clk_c), .Q(data_buffer_reg[395])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i395.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i396 (.D(data_buffer_reg_959__N_3020[396]), .SP(clk_c_enable_1000), 
            .CK(clk_c), .Q(data_buffer_reg[396])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i396.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i400 (.D(data_buffer_reg_959__N_3020[400]), .SP(clk_c_enable_1050), 
            .CK(clk_c), .Q(data_buffer_reg[400])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i400.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i401 (.D(data_buffer_reg_959__N_3020[401]), .SP(clk_c_enable_1050), 
            .CK(clk_c), .Q(data_buffer_reg[401])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i401.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i402 (.D(data_buffer_reg_959__N_3020[402]), .SP(clk_c_enable_1050), 
            .CK(clk_c), .Q(data_buffer_reg[402])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i402.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i403 (.D(data_buffer_reg_959__N_3020[403]), .SP(clk_c_enable_1050), 
            .CK(clk_c), .Q(data_buffer_reg[403])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i403.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i404 (.D(data_buffer_reg_959__N_3020[404]), .SP(clk_c_enable_1050), 
            .CK(clk_c), .Q(data_buffer_reg[404])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i404.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i408 (.D(data_buffer_reg_959__N_3020[408]), .SP(clk_c_enable_1050), 
            .CK(clk_c), .Q(data_buffer_reg[408])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i408.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i409 (.D(data_buffer_reg_959__N_3020[409]), .SP(clk_c_enable_1050), 
            .CK(clk_c), .Q(data_buffer_reg[409])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i409.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i410 (.D(data_buffer_reg_959__N_3020[410]), .SP(clk_c_enable_1050), 
            .CK(clk_c), .Q(data_buffer_reg[410])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i410.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i411 (.D(data_buffer_reg_959__N_3020[411]), .SP(clk_c_enable_1050), 
            .CK(clk_c), .Q(data_buffer_reg[411])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i411.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i412 (.D(data_buffer_reg_959__N_3020[412]), .SP(clk_c_enable_1050), 
            .CK(clk_c), .Q(data_buffer_reg[412])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i412.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i416 (.D(data_buffer_reg_959__N_3020[416]), .SP(clk_c_enable_1050), 
            .CK(clk_c), .Q(data_buffer_reg[416])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i416.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i417 (.D(data_buffer_reg_959__N_3020[417]), .SP(clk_c_enable_1050), 
            .CK(clk_c), .Q(data_buffer_reg[417])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i417.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i418 (.D(data_buffer_reg_959__N_3020[418]), .SP(clk_c_enable_1050), 
            .CK(clk_c), .Q(data_buffer_reg[418])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i418.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i419 (.D(data_buffer_reg_959__N_3020[419]), .SP(clk_c_enable_1050), 
            .CK(clk_c), .Q(data_buffer_reg[419])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i419.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i420 (.D(data_buffer_reg_959__N_3020[420]), .SP(clk_c_enable_1050), 
            .CK(clk_c), .Q(data_buffer_reg[420])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i420.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i424 (.D(data_buffer_reg_959__N_3020[424]), .SP(clk_c_enable_1050), 
            .CK(clk_c), .Q(data_buffer_reg[424])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i424.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i425 (.D(data_buffer_reg_959__N_3020[425]), .SP(clk_c_enable_1050), 
            .CK(clk_c), .Q(data_buffer_reg[425])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i425.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i426 (.D(data_buffer_reg_959__N_3020[426]), .SP(clk_c_enable_1050), 
            .CK(clk_c), .Q(data_buffer_reg[426])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i426.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i427 (.D(data_buffer_reg_959__N_3020[427]), .SP(clk_c_enable_1050), 
            .CK(clk_c), .Q(data_buffer_reg[427])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i427.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i428 (.D(data_buffer_reg_959__N_3020[428]), .SP(clk_c_enable_1050), 
            .CK(clk_c), .Q(data_buffer_reg[428])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i428.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i432 (.D(data_buffer_reg_959__N_3020[432]), .SP(clk_c_enable_1050), 
            .CK(clk_c), .Q(data_buffer_reg[432])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i432.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i433 (.D(data_buffer_reg_959__N_3020[433]), .SP(clk_c_enable_1050), 
            .CK(clk_c), .Q(data_buffer_reg[433])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i433.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i434 (.D(data_buffer_reg_959__N_3020[434]), .SP(clk_c_enable_1050), 
            .CK(clk_c), .Q(data_buffer_reg[434])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i434.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i435 (.D(data_buffer_reg_959__N_3020[435]), .SP(clk_c_enable_1050), 
            .CK(clk_c), .Q(data_buffer_reg[435])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i435.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i436 (.D(data_buffer_reg_959__N_3020[436]), .SP(clk_c_enable_1050), 
            .CK(clk_c), .Q(data_buffer_reg[436])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i436.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i440 (.D(data_buffer_reg_959__N_3020[440]), .SP(clk_c_enable_1050), 
            .CK(clk_c), .Q(data_buffer_reg[440])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i440.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i441 (.D(data_buffer_reg_959__N_3020[441]), .SP(clk_c_enable_1050), 
            .CK(clk_c), .Q(data_buffer_reg[441])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i441.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i442 (.D(data_buffer_reg_959__N_3020[442]), .SP(clk_c_enable_1050), 
            .CK(clk_c), .Q(data_buffer_reg[442])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i442.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i443 (.D(data_buffer_reg_959__N_3020[443]), .SP(clk_c_enable_1050), 
            .CK(clk_c), .Q(data_buffer_reg[443])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i443.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i444 (.D(data_buffer_reg_959__N_3020[444]), .SP(clk_c_enable_1050), 
            .CK(clk_c), .Q(data_buffer_reg[444])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i444.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i448 (.D(data_buffer_reg_959__N_3020[448]), .SP(clk_c_enable_1050), 
            .CK(clk_c), .Q(data_buffer_reg[448])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i448.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i449 (.D(data_buffer_reg_959__N_3020[449]), .SP(clk_c_enable_1050), 
            .CK(clk_c), .Q(data_buffer_reg[449])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i449.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i450 (.D(data_buffer_reg_959__N_3020[450]), .SP(clk_c_enable_1050), 
            .CK(clk_c), .Q(data_buffer_reg[450])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i450.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i451 (.D(data_buffer_reg_959__N_3020[451]), .SP(clk_c_enable_1050), 
            .CK(clk_c), .Q(data_buffer_reg[451])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i451.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i452 (.D(data_buffer_reg_959__N_3020[452]), .SP(clk_c_enable_1050), 
            .CK(clk_c), .Q(data_buffer_reg[452])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i452.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i456 (.D(data_buffer_reg_959__N_3020[456]), .SP(clk_c_enable_1050), 
            .CK(clk_c), .Q(data_buffer_reg[456])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i456.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i457 (.D(data_buffer_reg_959__N_3020[457]), .SP(clk_c_enable_1050), 
            .CK(clk_c), .Q(data_buffer_reg[457])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i457.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i458 (.D(data_buffer_reg_959__N_3020[458]), .SP(clk_c_enable_1050), 
            .CK(clk_c), .Q(data_buffer_reg[458])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i458.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i459 (.D(data_buffer_reg_959__N_3020[459]), .SP(clk_c_enable_1050), 
            .CK(clk_c), .Q(data_buffer_reg[459])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i459.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i460 (.D(data_buffer_reg_959__N_3020[460]), .SP(clk_c_enable_1050), 
            .CK(clk_c), .Q(data_buffer_reg[460])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i460.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i464 (.D(data_buffer_reg_959__N_3020[464]), .SP(clk_c_enable_1050), 
            .CK(clk_c), .Q(data_buffer_reg[464])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i464.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i465 (.D(data_buffer_reg_959__N_3020[465]), .SP(clk_c_enable_1050), 
            .CK(clk_c), .Q(data_buffer_reg[465])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i465.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i466 (.D(data_buffer_reg_959__N_3020[466]), .SP(clk_c_enable_1050), 
            .CK(clk_c), .Q(data_buffer_reg[466])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i466.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i467 (.D(data_buffer_reg_959__N_3020[467]), .SP(clk_c_enable_1050), 
            .CK(clk_c), .Q(data_buffer_reg[467])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i467.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i468 (.D(data_buffer_reg_959__N_3020[468]), .SP(clk_c_enable_1050), 
            .CK(clk_c), .Q(data_buffer_reg[468])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i468.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i472 (.D(data_buffer_reg_959__N_3020[472]), .SP(clk_c_enable_1050), 
            .CK(clk_c), .Q(data_buffer_reg[472])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i472.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i473 (.D(data_buffer_reg_959__N_3020[473]), .SP(clk_c_enable_1050), 
            .CK(clk_c), .Q(data_buffer_reg[473])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i473.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i474 (.D(data_buffer_reg_959__N_3020[474]), .SP(clk_c_enable_1050), 
            .CK(clk_c), .Q(data_buffer_reg[474])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i474.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i475 (.D(data_buffer_reg_959__N_3020[475]), .SP(clk_c_enable_1050), 
            .CK(clk_c), .Q(data_buffer_reg[475])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i475.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i476 (.D(data_buffer_reg_959__N_3020[476]), .SP(clk_c_enable_1050), 
            .CK(clk_c), .Q(data_buffer_reg[476])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i476.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i480 (.D(data_buffer_reg_959__N_3020[480]), .SP(clk_c_enable_1100), 
            .CK(clk_c), .Q(data_buffer_reg[480])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i480.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i481 (.D(data_buffer_reg_959__N_3020[481]), .SP(clk_c_enable_1100), 
            .CK(clk_c), .Q(data_buffer_reg[481])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i481.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i482 (.D(data_buffer_reg_959__N_3020[482]), .SP(clk_c_enable_1100), 
            .CK(clk_c), .Q(data_buffer_reg[482])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i482.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i483 (.D(data_buffer_reg_959__N_3020[483]), .SP(clk_c_enable_1100), 
            .CK(clk_c), .Q(data_buffer_reg[483])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i483.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i484 (.D(data_buffer_reg_959__N_3020[484]), .SP(clk_c_enable_1100), 
            .CK(clk_c), .Q(data_buffer_reg[484])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i484.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i488 (.D(data_buffer_reg_959__N_3020[488]), .SP(clk_c_enable_1100), 
            .CK(clk_c), .Q(data_buffer_reg[488])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i488.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i489 (.D(data_buffer_reg_959__N_3020[489]), .SP(clk_c_enable_1100), 
            .CK(clk_c), .Q(data_buffer_reg[489])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i489.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i490 (.D(data_buffer_reg_959__N_3020[490]), .SP(clk_c_enable_1100), 
            .CK(clk_c), .Q(data_buffer_reg[490])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i490.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i491 (.D(data_buffer_reg_959__N_3020[491]), .SP(clk_c_enable_1100), 
            .CK(clk_c), .Q(data_buffer_reg[491])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i491.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i492 (.D(data_buffer_reg_959__N_3020[492]), .SP(clk_c_enable_1100), 
            .CK(clk_c), .Q(data_buffer_reg[492])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i492.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i496 (.D(data_buffer_reg_959__N_3020[496]), .SP(clk_c_enable_1100), 
            .CK(clk_c), .Q(data_buffer_reg[496])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i496.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i497 (.D(data_buffer_reg_959__N_3020[497]), .SP(clk_c_enable_1100), 
            .CK(clk_c), .Q(data_buffer_reg[497])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i497.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i498 (.D(data_buffer_reg_959__N_3020[498]), .SP(clk_c_enable_1100), 
            .CK(clk_c), .Q(data_buffer_reg[498])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i498.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i499 (.D(data_buffer_reg_959__N_3020[499]), .SP(clk_c_enable_1100), 
            .CK(clk_c), .Q(data_buffer_reg[499])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i499.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i500 (.D(data_buffer_reg_959__N_3020[500]), .SP(clk_c_enable_1100), 
            .CK(clk_c), .Q(data_buffer_reg[500])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i500.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i504 (.D(data_buffer_reg_959__N_3020[504]), .SP(clk_c_enable_1100), 
            .CK(clk_c), .Q(data_buffer_reg[504])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i504.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i505 (.D(data_buffer_reg_959__N_3020[505]), .SP(clk_c_enable_1100), 
            .CK(clk_c), .Q(data_buffer_reg[505])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i505.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i506 (.D(data_buffer_reg_959__N_3020[506]), .SP(clk_c_enable_1100), 
            .CK(clk_c), .Q(data_buffer_reg[506])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i506.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i507 (.D(data_buffer_reg_959__N_3020[507]), .SP(clk_c_enable_1100), 
            .CK(clk_c), .Q(data_buffer_reg[507])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i507.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i508 (.D(data_buffer_reg_959__N_3020[508]), .SP(clk_c_enable_1100), 
            .CK(clk_c), .Q(data_buffer_reg[508])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i508.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i512 (.D(data_buffer_reg_959__N_3020[512]), .SP(clk_c_enable_1100), 
            .CK(clk_c), .Q(data_buffer_reg[512])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i512.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i513 (.D(data_buffer_reg_959__N_3020[513]), .SP(clk_c_enable_1100), 
            .CK(clk_c), .Q(data_buffer_reg[513])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i513.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i514 (.D(data_buffer_reg_959__N_3020[514]), .SP(clk_c_enable_1100), 
            .CK(clk_c), .Q(data_buffer_reg[514])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i514.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i515 (.D(data_buffer_reg_959__N_3020[515]), .SP(clk_c_enable_1100), 
            .CK(clk_c), .Q(data_buffer_reg[515])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i515.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i516 (.D(data_buffer_reg_959__N_3020[516]), .SP(clk_c_enable_1100), 
            .CK(clk_c), .Q(data_buffer_reg[516])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i516.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i520 (.D(data_buffer_reg_959__N_3020[520]), .SP(clk_c_enable_1100), 
            .CK(clk_c), .Q(data_buffer_reg[520])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i520.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i521 (.D(data_buffer_reg_959__N_3020[521]), .SP(clk_c_enable_1100), 
            .CK(clk_c), .Q(data_buffer_reg[521])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i521.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i522 (.D(data_buffer_reg_959__N_3020[522]), .SP(clk_c_enable_1100), 
            .CK(clk_c), .Q(data_buffer_reg[522])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i522.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i523 (.D(data_buffer_reg_959__N_3020[523]), .SP(clk_c_enable_1100), 
            .CK(clk_c), .Q(data_buffer_reg[523])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i523.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i524 (.D(data_buffer_reg_959__N_3020[524]), .SP(clk_c_enable_1100), 
            .CK(clk_c), .Q(data_buffer_reg[524])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i524.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i528 (.D(data_buffer_reg_959__N_3020[528]), .SP(clk_c_enable_1100), 
            .CK(clk_c), .Q(data_buffer_reg[528])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i528.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i529 (.D(data_buffer_reg_959__N_3020[529]), .SP(clk_c_enable_1100), 
            .CK(clk_c), .Q(data_buffer_reg[529])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i529.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i530 (.D(data_buffer_reg_959__N_3020[530]), .SP(clk_c_enable_1100), 
            .CK(clk_c), .Q(data_buffer_reg[530])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i530.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i531 (.D(data_buffer_reg_959__N_3020[531]), .SP(clk_c_enable_1100), 
            .CK(clk_c), .Q(data_buffer_reg[531])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i531.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i532 (.D(data_buffer_reg_959__N_3020[532]), .SP(clk_c_enable_1100), 
            .CK(clk_c), .Q(data_buffer_reg[532])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i532.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i536 (.D(data_buffer_reg_959__N_3020[536]), .SP(clk_c_enable_1100), 
            .CK(clk_c), .Q(data_buffer_reg[536])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i536.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i537 (.D(data_buffer_reg_959__N_3020[537]), .SP(clk_c_enable_1100), 
            .CK(clk_c), .Q(data_buffer_reg[537])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i537.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i538 (.D(data_buffer_reg_959__N_3020[538]), .SP(clk_c_enable_1100), 
            .CK(clk_c), .Q(data_buffer_reg[538])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i538.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i539 (.D(data_buffer_reg_959__N_3020[539]), .SP(clk_c_enable_1100), 
            .CK(clk_c), .Q(data_buffer_reg[539])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i539.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i540 (.D(data_buffer_reg_959__N_3020[540]), .SP(clk_c_enable_1100), 
            .CK(clk_c), .Q(data_buffer_reg[540])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i540.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i544 (.D(data_buffer_reg_959__N_3020[544]), .SP(clk_c_enable_1100), 
            .CK(clk_c), .Q(data_buffer_reg[544])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i544.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i545 (.D(data_buffer_reg_959__N_3020[545]), .SP(clk_c_enable_1100), 
            .CK(clk_c), .Q(data_buffer_reg[545])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i545.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i546 (.D(data_buffer_reg_959__N_3020[546]), .SP(clk_c_enable_1100), 
            .CK(clk_c), .Q(data_buffer_reg[546])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i546.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i547 (.D(data_buffer_reg_959__N_3020[547]), .SP(clk_c_enable_1100), 
            .CK(clk_c), .Q(data_buffer_reg[547])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i547.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i548 (.D(data_buffer_reg_959__N_3020[548]), .SP(clk_c_enable_1100), 
            .CK(clk_c), .Q(data_buffer_reg[548])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i548.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i552 (.D(data_buffer_reg_959__N_3020[552]), .SP(clk_c_enable_1100), 
            .CK(clk_c), .Q(data_buffer_reg[552])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i552.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i553 (.D(data_buffer_reg_959__N_3020[553]), .SP(clk_c_enable_1100), 
            .CK(clk_c), .Q(data_buffer_reg[553])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i553.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i554 (.D(data_buffer_reg_959__N_3020[554]), .SP(clk_c_enable_1100), 
            .CK(clk_c), .Q(data_buffer_reg[554])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i554.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i555 (.D(data_buffer_reg_959__N_3020[555]), .SP(clk_c_enable_1100), 
            .CK(clk_c), .Q(data_buffer_reg[555])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i555.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i556 (.D(data_buffer_reg_959__N_3020[556]), .SP(clk_c_enable_1100), 
            .CK(clk_c), .Q(data_buffer_reg[556])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i556.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i560 (.D(data_buffer_reg_959__N_3020[560]), .SP(clk_c_enable_1150), 
            .CK(clk_c), .Q(data_buffer_reg[560])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i560.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i561 (.D(data_buffer_reg_959__N_3020[561]), .SP(clk_c_enable_1150), 
            .CK(clk_c), .Q(data_buffer_reg[561])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i561.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i562 (.D(data_buffer_reg_959__N_3020[562]), .SP(clk_c_enable_1150), 
            .CK(clk_c), .Q(data_buffer_reg[562])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i562.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i563 (.D(data_buffer_reg_959__N_3020[563]), .SP(clk_c_enable_1150), 
            .CK(clk_c), .Q(data_buffer_reg[563])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i563.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i564 (.D(data_buffer_reg_959__N_3020[564]), .SP(clk_c_enable_1150), 
            .CK(clk_c), .Q(data_buffer_reg[564])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i564.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i568 (.D(data_buffer_reg_959__N_3020[568]), .SP(clk_c_enable_1150), 
            .CK(clk_c), .Q(data_buffer_reg[568])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i568.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i569 (.D(data_buffer_reg_959__N_3020[569]), .SP(clk_c_enable_1150), 
            .CK(clk_c), .Q(data_buffer_reg[569])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i569.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i570 (.D(data_buffer_reg_959__N_3020[570]), .SP(clk_c_enable_1150), 
            .CK(clk_c), .Q(data_buffer_reg[570])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i570.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i571 (.D(data_buffer_reg_959__N_3020[571]), .SP(clk_c_enable_1150), 
            .CK(clk_c), .Q(data_buffer_reg[571])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i571.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i572 (.D(data_buffer_reg_959__N_3020[572]), .SP(clk_c_enable_1150), 
            .CK(clk_c), .Q(data_buffer_reg[572])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i572.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i576 (.D(data_buffer_reg_959__N_3020[576]), .SP(clk_c_enable_1150), 
            .CK(clk_c), .Q(data_buffer_reg[576])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i576.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i577 (.D(data_buffer_reg_959__N_3020[577]), .SP(clk_c_enable_1150), 
            .CK(clk_c), .Q(data_buffer_reg[577])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i577.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i578 (.D(data_buffer_reg_959__N_3020[578]), .SP(clk_c_enable_1150), 
            .CK(clk_c), .Q(data_buffer_reg[578])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i578.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i579 (.D(data_buffer_reg_959__N_3020[579]), .SP(clk_c_enable_1150), 
            .CK(clk_c), .Q(data_buffer_reg[579])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i579.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i580 (.D(data_buffer_reg_959__N_3020[580]), .SP(clk_c_enable_1150), 
            .CK(clk_c), .Q(data_buffer_reg[580])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i580.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i584 (.D(data_buffer_reg_959__N_3020[584]), .SP(clk_c_enable_1150), 
            .CK(clk_c), .Q(data_buffer_reg[584])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i584.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i585 (.D(data_buffer_reg_959__N_3020[585]), .SP(clk_c_enable_1150), 
            .CK(clk_c), .Q(data_buffer_reg[585])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i585.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i586 (.D(data_buffer_reg_959__N_3020[586]), .SP(clk_c_enable_1150), 
            .CK(clk_c), .Q(data_buffer_reg[586])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i586.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i587 (.D(data_buffer_reg_959__N_3020[587]), .SP(clk_c_enable_1150), 
            .CK(clk_c), .Q(data_buffer_reg[587])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i587.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i588 (.D(data_buffer_reg_959__N_3020[588]), .SP(clk_c_enable_1150), 
            .CK(clk_c), .Q(data_buffer_reg[588])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i588.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i592 (.D(data_buffer_reg_959__N_3020[592]), .SP(clk_c_enable_1150), 
            .CK(clk_c), .Q(data_buffer_reg[592])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i592.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i593 (.D(data_buffer_reg_959__N_3020[593]), .SP(clk_c_enable_1150), 
            .CK(clk_c), .Q(data_buffer_reg[593])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i593.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i594 (.D(data_buffer_reg_959__N_3020[594]), .SP(clk_c_enable_1150), 
            .CK(clk_c), .Q(data_buffer_reg[594])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i594.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i595 (.D(data_buffer_reg_959__N_3020[595]), .SP(clk_c_enable_1150), 
            .CK(clk_c), .Q(data_buffer_reg[595])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i595.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i596 (.D(data_buffer_reg_959__N_3020[596]), .SP(clk_c_enable_1150), 
            .CK(clk_c), .Q(data_buffer_reg[596])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i596.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i600 (.D(data_buffer_reg_959__N_3020[600]), .SP(clk_c_enable_1150), 
            .CK(clk_c), .Q(data_buffer_reg[600])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i600.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i601 (.D(data_buffer_reg_959__N_3020[601]), .SP(clk_c_enable_1150), 
            .CK(clk_c), .Q(data_buffer_reg[601])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i601.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i602 (.D(data_buffer_reg_959__N_3020[602]), .SP(clk_c_enable_1150), 
            .CK(clk_c), .Q(data_buffer_reg[602])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i602.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i603 (.D(data_buffer_reg_959__N_3020[603]), .SP(clk_c_enable_1150), 
            .CK(clk_c), .Q(data_buffer_reg[603])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i603.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i604 (.D(data_buffer_reg_959__N_3020[604]), .SP(clk_c_enable_1150), 
            .CK(clk_c), .Q(data_buffer_reg[604])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i604.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i608 (.D(data_buffer_reg_959__N_3020[608]), .SP(clk_c_enable_1150), 
            .CK(clk_c), .Q(data_buffer_reg[608])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i608.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i609 (.D(data_buffer_reg_959__N_3020[609]), .SP(clk_c_enable_1150), 
            .CK(clk_c), .Q(data_buffer_reg[609])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i609.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i610 (.D(data_buffer_reg_959__N_3020[610]), .SP(clk_c_enable_1150), 
            .CK(clk_c), .Q(data_buffer_reg[610])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i610.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i611 (.D(data_buffer_reg_959__N_3020[611]), .SP(clk_c_enable_1150), 
            .CK(clk_c), .Q(data_buffer_reg[611])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i611.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i612 (.D(data_buffer_reg_959__N_3020[612]), .SP(clk_c_enable_1150), 
            .CK(clk_c), .Q(data_buffer_reg[612])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i612.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i616 (.D(data_buffer_reg_959__N_3020[616]), .SP(clk_c_enable_1150), 
            .CK(clk_c), .Q(data_buffer_reg[616])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i616.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i617 (.D(data_buffer_reg_959__N_3020[617]), .SP(clk_c_enable_1150), 
            .CK(clk_c), .Q(data_buffer_reg[617])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i617.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i618 (.D(data_buffer_reg_959__N_3020[618]), .SP(clk_c_enable_1150), 
            .CK(clk_c), .Q(data_buffer_reg[618])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i618.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i619 (.D(data_buffer_reg_959__N_3020[619]), .SP(clk_c_enable_1150), 
            .CK(clk_c), .Q(data_buffer_reg[619])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i619.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i620 (.D(data_buffer_reg_959__N_3020[620]), .SP(clk_c_enable_1150), 
            .CK(clk_c), .Q(data_buffer_reg[620])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i620.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i624 (.D(data_buffer_reg_959__N_3020[624]), .SP(clk_c_enable_1150), 
            .CK(clk_c), .Q(data_buffer_reg[624])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i624.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i625 (.D(data_buffer_reg_959__N_3020[625]), .SP(clk_c_enable_1150), 
            .CK(clk_c), .Q(data_buffer_reg[625])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i625.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i626 (.D(data_buffer_reg_959__N_3020[626]), .SP(clk_c_enable_1150), 
            .CK(clk_c), .Q(data_buffer_reg[626])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i626.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i627 (.D(data_buffer_reg_959__N_3020[627]), .SP(clk_c_enable_1150), 
            .CK(clk_c), .Q(data_buffer_reg[627])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i627.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i628 (.D(data_buffer_reg_959__N_3020[628]), .SP(clk_c_enable_1150), 
            .CK(clk_c), .Q(data_buffer_reg[628])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i628.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i632 (.D(data_buffer_reg_959__N_3020[632]), .SP(clk_c_enable_1150), 
            .CK(clk_c), .Q(data_buffer_reg[632])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i632.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i633 (.D(data_buffer_reg_959__N_3020[633]), .SP(clk_c_enable_1150), 
            .CK(clk_c), .Q(data_buffer_reg[633])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i633.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i634 (.D(data_buffer_reg_959__N_3020[634]), .SP(clk_c_enable_1150), 
            .CK(clk_c), .Q(data_buffer_reg[634])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i634.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i635 (.D(data_buffer_reg_959__N_3020[635]), .SP(clk_c_enable_1150), 
            .CK(clk_c), .Q(data_buffer_reg[635])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i635.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i636 (.D(data_buffer_reg_959__N_3020[636]), .SP(clk_c_enable_1150), 
            .CK(clk_c), .Q(data_buffer_reg[636])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i636.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i640 (.D(data_buffer_reg_959__N_3020[640]), .SP(clk_c_enable_1200), 
            .CK(clk_c), .Q(data_buffer_reg[640])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i640.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i641 (.D(data_buffer_reg_959__N_3020[641]), .SP(clk_c_enable_1200), 
            .CK(clk_c), .Q(data_buffer_reg[641])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i641.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i642 (.D(data_buffer_reg_959__N_3020[642]), .SP(clk_c_enable_1200), 
            .CK(clk_c), .Q(data_buffer_reg[642])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i642.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i643 (.D(data_buffer_reg_959__N_3020[643]), .SP(clk_c_enable_1200), 
            .CK(clk_c), .Q(data_buffer_reg[643])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i643.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i644 (.D(data_buffer_reg_959__N_3020[644]), .SP(clk_c_enable_1200), 
            .CK(clk_c), .Q(data_buffer_reg[644])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i644.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i648 (.D(data_buffer_reg_959__N_3020[648]), .SP(clk_c_enable_1200), 
            .CK(clk_c), .Q(data_buffer_reg[648])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i648.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i649 (.D(data_buffer_reg_959__N_3020[649]), .SP(clk_c_enable_1200), 
            .CK(clk_c), .Q(data_buffer_reg[649])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i649.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i650 (.D(data_buffer_reg_959__N_3020[650]), .SP(clk_c_enable_1200), 
            .CK(clk_c), .Q(data_buffer_reg[650])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i650.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i651 (.D(data_buffer_reg_959__N_3020[651]), .SP(clk_c_enable_1200), 
            .CK(clk_c), .Q(data_buffer_reg[651])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i651.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i652 (.D(data_buffer_reg_959__N_3020[652]), .SP(clk_c_enable_1200), 
            .CK(clk_c), .Q(data_buffer_reg[652])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i652.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i656 (.D(data_buffer_reg_959__N_3020[656]), .SP(clk_c_enable_1200), 
            .CK(clk_c), .Q(data_buffer_reg[656])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i656.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i657 (.D(data_buffer_reg_959__N_3020[657]), .SP(clk_c_enable_1200), 
            .CK(clk_c), .Q(data_buffer_reg[657])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i657.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i658 (.D(data_buffer_reg_959__N_3020[658]), .SP(clk_c_enable_1200), 
            .CK(clk_c), .Q(data_buffer_reg[658])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i658.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i659 (.D(data_buffer_reg_959__N_3020[659]), .SP(clk_c_enable_1200), 
            .CK(clk_c), .Q(data_buffer_reg[659])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i659.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i660 (.D(data_buffer_reg_959__N_3020[660]), .SP(clk_c_enable_1200), 
            .CK(clk_c), .Q(data_buffer_reg[660])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i660.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i664 (.D(data_buffer_reg_959__N_3020[664]), .SP(clk_c_enable_1200), 
            .CK(clk_c), .Q(data_buffer_reg[664])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i664.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i665 (.D(data_buffer_reg_959__N_3020[665]), .SP(clk_c_enable_1200), 
            .CK(clk_c), .Q(data_buffer_reg[665])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i665.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i666 (.D(data_buffer_reg_959__N_3020[666]), .SP(clk_c_enable_1200), 
            .CK(clk_c), .Q(data_buffer_reg[666])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i666.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i667 (.D(data_buffer_reg_959__N_3020[667]), .SP(clk_c_enable_1200), 
            .CK(clk_c), .Q(data_buffer_reg[667])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i667.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i668 (.D(data_buffer_reg_959__N_3020[668]), .SP(clk_c_enable_1200), 
            .CK(clk_c), .Q(data_buffer_reg[668])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i668.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i672 (.D(data_buffer_reg_959__N_3020[672]), .SP(clk_c_enable_1200), 
            .CK(clk_c), .Q(data_buffer_reg[672])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i672.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i673 (.D(data_buffer_reg_959__N_3020[673]), .SP(clk_c_enable_1200), 
            .CK(clk_c), .Q(data_buffer_reg[673])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i673.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i674 (.D(data_buffer_reg_959__N_3020[674]), .SP(clk_c_enable_1200), 
            .CK(clk_c), .Q(data_buffer_reg[674])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i674.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i675 (.D(data_buffer_reg_959__N_3020[675]), .SP(clk_c_enable_1200), 
            .CK(clk_c), .Q(data_buffer_reg[675])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i675.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i676 (.D(data_buffer_reg_959__N_3020[676]), .SP(clk_c_enable_1200), 
            .CK(clk_c), .Q(data_buffer_reg[676])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i676.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i680 (.D(data_buffer_reg_959__N_3020[680]), .SP(clk_c_enable_1200), 
            .CK(clk_c), .Q(data_buffer_reg[680])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i680.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i681 (.D(data_buffer_reg_959__N_3020[681]), .SP(clk_c_enable_1200), 
            .CK(clk_c), .Q(data_buffer_reg[681])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i681.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i682 (.D(data_buffer_reg_959__N_3020[682]), .SP(clk_c_enable_1200), 
            .CK(clk_c), .Q(data_buffer_reg[682])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i682.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i683 (.D(data_buffer_reg_959__N_3020[683]), .SP(clk_c_enable_1200), 
            .CK(clk_c), .Q(data_buffer_reg[683])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i683.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i684 (.D(data_buffer_reg_959__N_3020[684]), .SP(clk_c_enable_1200), 
            .CK(clk_c), .Q(data_buffer_reg[684])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i684.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i688 (.D(data_buffer_reg_959__N_3020[688]), .SP(clk_c_enable_1200), 
            .CK(clk_c), .Q(data_buffer_reg[688])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i688.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i689 (.D(data_buffer_reg_959__N_3020[689]), .SP(clk_c_enable_1200), 
            .CK(clk_c), .Q(data_buffer_reg[689])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i689.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i690 (.D(data_buffer_reg_959__N_3020[690]), .SP(clk_c_enable_1200), 
            .CK(clk_c), .Q(data_buffer_reg[690])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i690.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i691 (.D(data_buffer_reg_959__N_3020[691]), .SP(clk_c_enable_1200), 
            .CK(clk_c), .Q(data_buffer_reg[691])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i691.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i692 (.D(data_buffer_reg_959__N_3020[692]), .SP(clk_c_enable_1200), 
            .CK(clk_c), .Q(data_buffer_reg[692])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i692.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i696 (.D(data_buffer_reg_959__N_3020[696]), .SP(clk_c_enable_1200), 
            .CK(clk_c), .Q(data_buffer_reg[696])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i696.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i697 (.D(data_buffer_reg_959__N_3020[697]), .SP(clk_c_enable_1200), 
            .CK(clk_c), .Q(data_buffer_reg[697])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i697.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i698 (.D(data_buffer_reg_959__N_3020[698]), .SP(clk_c_enable_1200), 
            .CK(clk_c), .Q(data_buffer_reg[698])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i698.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i699 (.D(data_buffer_reg_959__N_3020[699]), .SP(clk_c_enable_1200), 
            .CK(clk_c), .Q(data_buffer_reg[699])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i699.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i700 (.D(data_buffer_reg_959__N_3020[700]), .SP(clk_c_enable_1200), 
            .CK(clk_c), .Q(data_buffer_reg[700])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i700.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i704 (.D(data_buffer_reg_959__N_3020[704]), .SP(clk_c_enable_1200), 
            .CK(clk_c), .Q(data_buffer_reg[704])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i704.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i705 (.D(data_buffer_reg_959__N_3020[705]), .SP(clk_c_enable_1200), 
            .CK(clk_c), .Q(data_buffer_reg[705])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i705.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i706 (.D(data_buffer_reg_959__N_3020[706]), .SP(clk_c_enable_1200), 
            .CK(clk_c), .Q(data_buffer_reg[706])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i706.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i707 (.D(data_buffer_reg_959__N_3020[707]), .SP(clk_c_enable_1200), 
            .CK(clk_c), .Q(data_buffer_reg[707])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i707.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i708 (.D(data_buffer_reg_959__N_3020[708]), .SP(clk_c_enable_1200), 
            .CK(clk_c), .Q(data_buffer_reg[708])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i708.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i712 (.D(data_buffer_reg_959__N_3020[712]), .SP(clk_c_enable_1200), 
            .CK(clk_c), .Q(data_buffer_reg[712])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i712.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i713 (.D(data_buffer_reg_959__N_3020[713]), .SP(clk_c_enable_1200), 
            .CK(clk_c), .Q(data_buffer_reg[713])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i713.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i714 (.D(data_buffer_reg_959__N_3020[714]), .SP(clk_c_enable_1200), 
            .CK(clk_c), .Q(data_buffer_reg[714])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i714.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i715 (.D(data_buffer_reg_959__N_3020[715]), .SP(clk_c_enable_1200), 
            .CK(clk_c), .Q(data_buffer_reg[715])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i715.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i716 (.D(data_buffer_reg_959__N_3020[716]), .SP(clk_c_enable_1200), 
            .CK(clk_c), .Q(data_buffer_reg[716])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i716.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i720 (.D(data_buffer_reg_959__N_3020[720]), .SP(clk_c_enable_1250), 
            .CK(clk_c), .Q(data_buffer_reg[720])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i720.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i721 (.D(data_buffer_reg_959__N_3020[721]), .SP(clk_c_enable_1250), 
            .CK(clk_c), .Q(data_buffer_reg[721])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i721.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i722 (.D(data_buffer_reg_959__N_3020[722]), .SP(clk_c_enable_1250), 
            .CK(clk_c), .Q(data_buffer_reg[722])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i722.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i723 (.D(data_buffer_reg_959__N_3020[723]), .SP(clk_c_enable_1250), 
            .CK(clk_c), .Q(data_buffer_reg[723])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i723.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i724 (.D(data_buffer_reg_959__N_3020[724]), .SP(clk_c_enable_1250), 
            .CK(clk_c), .Q(data_buffer_reg[724])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i724.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i728 (.D(data_buffer_reg_959__N_3020[728]), .SP(clk_c_enable_1250), 
            .CK(clk_c), .Q(data_buffer_reg[728])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i728.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i729 (.D(data_buffer_reg_959__N_3020[729]), .SP(clk_c_enable_1250), 
            .CK(clk_c), .Q(data_buffer_reg[729])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i729.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i730 (.D(data_buffer_reg_959__N_3020[730]), .SP(clk_c_enable_1250), 
            .CK(clk_c), .Q(data_buffer_reg[730])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i730.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i731 (.D(data_buffer_reg_959__N_3020[731]), .SP(clk_c_enable_1250), 
            .CK(clk_c), .Q(data_buffer_reg[731])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i731.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i732 (.D(data_buffer_reg_959__N_3020[732]), .SP(clk_c_enable_1250), 
            .CK(clk_c), .Q(data_buffer_reg[732])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i732.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i736 (.D(data_buffer_reg_959__N_3020[736]), .SP(clk_c_enable_1250), 
            .CK(clk_c), .Q(data_buffer_reg[736])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i736.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i737 (.D(data_buffer_reg_959__N_3020[737]), .SP(clk_c_enable_1250), 
            .CK(clk_c), .Q(data_buffer_reg[737])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i737.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i738 (.D(data_buffer_reg_959__N_3020[738]), .SP(clk_c_enable_1250), 
            .CK(clk_c), .Q(data_buffer_reg[738])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i738.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i739 (.D(data_buffer_reg_959__N_3020[739]), .SP(clk_c_enable_1250), 
            .CK(clk_c), .Q(data_buffer_reg[739])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i739.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i740 (.D(data_buffer_reg_959__N_3020[740]), .SP(clk_c_enable_1250), 
            .CK(clk_c), .Q(data_buffer_reg[740])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i740.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i744 (.D(data_buffer_reg_959__N_3020[744]), .SP(clk_c_enable_1250), 
            .CK(clk_c), .Q(data_buffer_reg[744])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i744.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i745 (.D(data_buffer_reg_959__N_3020[745]), .SP(clk_c_enable_1250), 
            .CK(clk_c), .Q(data_buffer_reg[745])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i745.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i746 (.D(data_buffer_reg_959__N_3020[746]), .SP(clk_c_enable_1250), 
            .CK(clk_c), .Q(data_buffer_reg[746])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i746.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i747 (.D(data_buffer_reg_959__N_3020[747]), .SP(clk_c_enable_1250), 
            .CK(clk_c), .Q(data_buffer_reg[747])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i747.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i748 (.D(data_buffer_reg_959__N_3020[748]), .SP(clk_c_enable_1250), 
            .CK(clk_c), .Q(data_buffer_reg[748])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i748.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i752 (.D(data_buffer_reg_959__N_3020[752]), .SP(clk_c_enable_1250), 
            .CK(clk_c), .Q(data_buffer_reg[752])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i752.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i753 (.D(data_buffer_reg_959__N_3020[753]), .SP(clk_c_enable_1250), 
            .CK(clk_c), .Q(data_buffer_reg[753])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i753.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i754 (.D(data_buffer_reg_959__N_3020[754]), .SP(clk_c_enable_1250), 
            .CK(clk_c), .Q(data_buffer_reg[754])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i754.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i755 (.D(data_buffer_reg_959__N_3020[755]), .SP(clk_c_enable_1250), 
            .CK(clk_c), .Q(data_buffer_reg[755])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i755.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i756 (.D(data_buffer_reg_959__N_3020[756]), .SP(clk_c_enable_1250), 
            .CK(clk_c), .Q(data_buffer_reg[756])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i756.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i760 (.D(data_buffer_reg_959__N_3020[760]), .SP(clk_c_enable_1250), 
            .CK(clk_c), .Q(data_buffer_reg[760])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i760.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i761 (.D(data_buffer_reg_959__N_3020[761]), .SP(clk_c_enable_1250), 
            .CK(clk_c), .Q(data_buffer_reg[761])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i761.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i762 (.D(data_buffer_reg_959__N_3020[762]), .SP(clk_c_enable_1250), 
            .CK(clk_c), .Q(data_buffer_reg[762])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i762.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i763 (.D(data_buffer_reg_959__N_3020[763]), .SP(clk_c_enable_1250), 
            .CK(clk_c), .Q(data_buffer_reg[763])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i763.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i764 (.D(data_buffer_reg_959__N_3020[764]), .SP(clk_c_enable_1250), 
            .CK(clk_c), .Q(data_buffer_reg[764])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i764.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i768 (.D(data_buffer_reg_959__N_3020[768]), .SP(clk_c_enable_1250), 
            .CK(clk_c), .Q(data_buffer_reg[768])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i768.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i769 (.D(data_buffer_reg_959__N_3020[769]), .SP(clk_c_enable_1250), 
            .CK(clk_c), .Q(data_buffer_reg[769])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i769.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i770 (.D(data_buffer_reg_959__N_3020[770]), .SP(clk_c_enable_1250), 
            .CK(clk_c), .Q(data_buffer_reg[770])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i770.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i771 (.D(data_buffer_reg_959__N_3020[771]), .SP(clk_c_enable_1250), 
            .CK(clk_c), .Q(data_buffer_reg[771])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i771.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i772 (.D(data_buffer_reg_959__N_3020[772]), .SP(clk_c_enable_1250), 
            .CK(clk_c), .Q(data_buffer_reg[772])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i772.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i776 (.D(data_buffer_reg_959__N_3020[776]), .SP(clk_c_enable_1250), 
            .CK(clk_c), .Q(data_buffer_reg[776])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i776.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i777 (.D(data_buffer_reg_959__N_3020[777]), .SP(clk_c_enable_1250), 
            .CK(clk_c), .Q(data_buffer_reg[777])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i777.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i778 (.D(data_buffer_reg_959__N_3020[778]), .SP(clk_c_enable_1250), 
            .CK(clk_c), .Q(data_buffer_reg[778])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i778.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i779 (.D(data_buffer_reg_959__N_3020[779]), .SP(clk_c_enable_1250), 
            .CK(clk_c), .Q(data_buffer_reg[779])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i779.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i780 (.D(data_buffer_reg_959__N_3020[780]), .SP(clk_c_enable_1250), 
            .CK(clk_c), .Q(data_buffer_reg[780])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i780.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i784 (.D(data_buffer_reg_959__N_3020[784]), .SP(clk_c_enable_1250), 
            .CK(clk_c), .Q(data_buffer_reg[784])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i784.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i785 (.D(data_buffer_reg_959__N_3020[785]), .SP(clk_c_enable_1250), 
            .CK(clk_c), .Q(data_buffer_reg[785])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i785.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i786 (.D(data_buffer_reg_959__N_3020[786]), .SP(clk_c_enable_1250), 
            .CK(clk_c), .Q(data_buffer_reg[786])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i786.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i787 (.D(data_buffer_reg_959__N_3020[787]), .SP(clk_c_enable_1250), 
            .CK(clk_c), .Q(data_buffer_reg[787])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i787.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i788 (.D(data_buffer_reg_959__N_3020[788]), .SP(clk_c_enable_1250), 
            .CK(clk_c), .Q(data_buffer_reg[788])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i788.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i792 (.D(data_buffer_reg_959__N_3020[792]), .SP(clk_c_enable_1250), 
            .CK(clk_c), .Q(data_buffer_reg[792])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i792.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i793 (.D(data_buffer_reg_959__N_3020[793]), .SP(clk_c_enable_1250), 
            .CK(clk_c), .Q(data_buffer_reg[793])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i793.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i794 (.D(data_buffer_reg_959__N_3020[794]), .SP(clk_c_enable_1250), 
            .CK(clk_c), .Q(data_buffer_reg[794])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i794.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i795 (.D(data_buffer_reg_959__N_3020[795]), .SP(clk_c_enable_1250), 
            .CK(clk_c), .Q(data_buffer_reg[795])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i795.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i796 (.D(data_buffer_reg_959__N_3020[796]), .SP(clk_c_enable_1250), 
            .CK(clk_c), .Q(data_buffer_reg[796])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i796.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i800 (.D(data_buffer_reg_959__N_3020[800]), .SP(clk_c_enable_1304), 
            .CK(clk_c), .Q(data_buffer_reg[800])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i800.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i801 (.D(data_buffer_reg_959__N_3020[801]), .SP(clk_c_enable_1304), 
            .CK(clk_c), .Q(data_buffer_reg[801])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i801.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i802 (.D(data_buffer_reg_959__N_3020[802]), .SP(clk_c_enable_1304), 
            .CK(clk_c), .Q(data_buffer_reg[802])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i802.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i803 (.D(data_buffer_reg_959__N_3020[803]), .SP(clk_c_enable_1304), 
            .CK(clk_c), .Q(data_buffer_reg[803])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i803.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i804 (.D(data_buffer_reg_959__N_3020[804]), .SP(clk_c_enable_1304), 
            .CK(clk_c), .Q(data_buffer_reg[804])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i804.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i808 (.D(data_buffer_reg_959__N_3020[808]), .SP(clk_c_enable_1304), 
            .CK(clk_c), .Q(data_buffer_reg[808])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i808.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i809 (.D(data_buffer_reg_959__N_3020[809]), .SP(clk_c_enable_1304), 
            .CK(clk_c), .Q(data_buffer_reg[809])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i809.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i810 (.D(data_buffer_reg_959__N_3020[810]), .SP(clk_c_enable_1304), 
            .CK(clk_c), .Q(data_buffer_reg[810])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i810.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i811 (.D(data_buffer_reg_959__N_3020[811]), .SP(clk_c_enable_1304), 
            .CK(clk_c), .Q(data_buffer_reg[811])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i811.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i812 (.D(data_buffer_reg_959__N_3020[812]), .SP(clk_c_enable_1304), 
            .CK(clk_c), .Q(data_buffer_reg[812])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i812.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i816 (.D(data_buffer_reg_959__N_3020[816]), .SP(clk_c_enable_1304), 
            .CK(clk_c), .Q(data_buffer_reg[816])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i816.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i817 (.D(data_buffer_reg_959__N_3020[817]), .SP(clk_c_enable_1304), 
            .CK(clk_c), .Q(data_buffer_reg[817])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i817.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i818 (.D(data_buffer_reg_959__N_3020[818]), .SP(clk_c_enable_1304), 
            .CK(clk_c), .Q(data_buffer_reg[818])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i818.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i819 (.D(data_buffer_reg_959__N_3020[819]), .SP(clk_c_enable_1304), 
            .CK(clk_c), .Q(data_buffer_reg[819])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i819.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i820 (.D(data_buffer_reg_959__N_3020[820]), .SP(clk_c_enable_1304), 
            .CK(clk_c), .Q(data_buffer_reg[820])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i820.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i824 (.D(data_buffer_reg_959__N_3020[824]), .SP(clk_c_enable_1304), 
            .CK(clk_c), .Q(data_buffer_reg[824])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i824.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i825 (.D(data_buffer_reg_959__N_3020[825]), .SP(clk_c_enable_1304), 
            .CK(clk_c), .Q(data_buffer_reg[825])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i825.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i826 (.D(data_buffer_reg_959__N_3020[826]), .SP(clk_c_enable_1304), 
            .CK(clk_c), .Q(data_buffer_reg[826])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i826.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i827 (.D(data_buffer_reg_959__N_3020[827]), .SP(clk_c_enable_1304), 
            .CK(clk_c), .Q(data_buffer_reg[827])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i827.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i828 (.D(data_buffer_reg_959__N_3020[828]), .SP(clk_c_enable_1304), 
            .CK(clk_c), .Q(data_buffer_reg[828])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i828.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i832 (.D(data_buffer_reg_959__N_3020[832]), .SP(clk_c_enable_1304), 
            .CK(clk_c), .Q(data_buffer_reg[832])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i832.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i833 (.D(data_buffer_reg_959__N_3020[833]), .SP(clk_c_enable_1304), 
            .CK(clk_c), .Q(data_buffer_reg[833])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i833.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i834 (.D(data_buffer_reg_959__N_3020[834]), .SP(clk_c_enable_1304), 
            .CK(clk_c), .Q(data_buffer_reg[834])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i834.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i835 (.D(data_buffer_reg_959__N_3020[835]), .SP(clk_c_enable_1304), 
            .CK(clk_c), .Q(data_buffer_reg[835])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i835.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i836 (.D(data_buffer_reg_959__N_3020[836]), .SP(clk_c_enable_1304), 
            .CK(clk_c), .Q(data_buffer_reg[836])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i836.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i840 (.D(data_buffer_reg_959__N_3020[840]), .SP(clk_c_enable_1304), 
            .CK(clk_c), .Q(data_buffer_reg[840])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i840.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i841 (.D(data_buffer_reg_959__N_3020[841]), .SP(clk_c_enable_1304), 
            .CK(clk_c), .Q(data_buffer_reg[841])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i841.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i842 (.D(data_buffer_reg_959__N_3020[842]), .SP(clk_c_enable_1304), 
            .CK(clk_c), .Q(data_buffer_reg[842])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i842.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i843 (.D(data_buffer_reg_959__N_3020[843]), .SP(clk_c_enable_1304), 
            .CK(clk_c), .Q(data_buffer_reg[843])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i843.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i844 (.D(data_buffer_reg_959__N_3020[844]), .SP(clk_c_enable_1304), 
            .CK(clk_c), .Q(data_buffer_reg[844])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i844.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i848 (.D(data_buffer_reg_959__N_3020[848]), .SP(clk_c_enable_1304), 
            .CK(clk_c), .Q(data_buffer_reg[848])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i848.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i849 (.D(data_buffer_reg_959__N_3020[849]), .SP(clk_c_enable_1304), 
            .CK(clk_c), .Q(data_buffer_reg[849])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i849.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i850 (.D(data_buffer_reg_959__N_3020[850]), .SP(clk_c_enable_1304), 
            .CK(clk_c), .Q(data_buffer_reg[850])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i850.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i851 (.D(data_buffer_reg_959__N_3020[851]), .SP(clk_c_enable_1304), 
            .CK(clk_c), .Q(data_buffer_reg[851])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i851.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i852 (.D(data_buffer_reg_959__N_3020[852]), .SP(clk_c_enable_1304), 
            .CK(clk_c), .Q(data_buffer_reg[852])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i852.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i856 (.D(data_buffer_reg_959__N_3020[856]), .SP(clk_c_enable_1304), 
            .CK(clk_c), .Q(data_buffer_reg[856])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i856.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i857 (.D(data_buffer_reg_959__N_3020[857]), .SP(clk_c_enable_1304), 
            .CK(clk_c), .Q(data_buffer_reg[857])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i857.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i858 (.D(data_buffer_reg_959__N_3020[858]), .SP(clk_c_enable_1304), 
            .CK(clk_c), .Q(data_buffer_reg[858])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i858.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i859 (.D(data_buffer_reg_959__N_3020[859]), .SP(clk_c_enable_1304), 
            .CK(clk_c), .Q(data_buffer_reg[859])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i859.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i860 (.D(data_buffer_reg_959__N_3020[860]), .SP(clk_c_enable_1304), 
            .CK(clk_c), .Q(data_buffer_reg[860])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i860.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i864 (.D(data_buffer_reg_959__N_3020[864]), .SP(clk_c_enable_1304), 
            .CK(clk_c), .Q(data_buffer_reg[864])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i864.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i865 (.D(data_buffer_reg_959__N_3020[865]), .SP(clk_c_enable_1304), 
            .CK(clk_c), .Q(data_buffer_reg[865])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i865.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i866 (.D(data_buffer_reg_959__N_3020[866]), .SP(clk_c_enable_1304), 
            .CK(clk_c), .Q(data_buffer_reg[866])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i866.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i867 (.D(data_buffer_reg_959__N_3020[867]), .SP(clk_c_enable_1304), 
            .CK(clk_c), .Q(data_buffer_reg[867])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i867.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i868 (.D(data_buffer_reg_959__N_3020[868]), .SP(clk_c_enable_1304), 
            .CK(clk_c), .Q(data_buffer_reg[868])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i868.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i872 (.D(data_buffer_reg_959__N_3020[872]), .SP(clk_c_enable_1304), 
            .CK(clk_c), .Q(data_buffer_reg[872])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i872.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i873 (.D(data_buffer_reg_959__N_3020[873]), .SP(clk_c_enable_1304), 
            .CK(clk_c), .Q(data_buffer_reg[873])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i873.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i874 (.D(data_buffer_reg_959__N_3020[874]), .SP(clk_c_enable_1304), 
            .CK(clk_c), .Q(data_buffer_reg[874])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i874.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i875 (.D(data_buffer_reg_959__N_3020[875]), .SP(clk_c_enable_1304), 
            .CK(clk_c), .Q(data_buffer_reg[875])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i875.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i876 (.D(data_buffer_reg_959__N_3020[876]), .SP(clk_c_enable_1304), 
            .CK(clk_c), .Q(data_buffer_reg[876])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i876.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i880 (.D(data_buffer_reg_959__N_3020[880]), .SP(clk_c_enable_1414), 
            .CK(clk_c), .Q(data_buffer_reg[880])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i880.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i881 (.D(data_buffer_reg_959__N_3020[881]), .SP(clk_c_enable_1414), 
            .CK(clk_c), .Q(data_buffer_reg[881])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i881.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i882 (.D(data_buffer_reg_959__N_3020[882]), .SP(clk_c_enable_1414), 
            .CK(clk_c), .Q(data_buffer_reg[882])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i882.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i883 (.D(data_buffer_reg_959__N_3020[883]), .SP(clk_c_enable_1414), 
            .CK(clk_c), .Q(data_buffer_reg[883])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i883.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i884 (.D(data_buffer_reg_959__N_3020[884]), .SP(clk_c_enable_1414), 
            .CK(clk_c), .Q(data_buffer_reg[884])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i884.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i888 (.D(data_buffer_reg_959__N_3020[888]), .SP(clk_c_enable_1414), 
            .CK(clk_c), .Q(data_buffer_reg[888])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i888.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i889 (.D(data_buffer_reg_959__N_3020[889]), .SP(clk_c_enable_1414), 
            .CK(clk_c), .Q(data_buffer_reg[889])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i889.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i890 (.D(data_buffer_reg_959__N_3020[890]), .SP(clk_c_enable_1414), 
            .CK(clk_c), .Q(data_buffer_reg[890])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i890.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i891 (.D(data_buffer_reg_959__N_3020[891]), .SP(clk_c_enable_1414), 
            .CK(clk_c), .Q(data_buffer_reg[891])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i891.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i892 (.D(data_buffer_reg_959__N_3020[892]), .SP(clk_c_enable_1414), 
            .CK(clk_c), .Q(data_buffer_reg[892])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i892.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i896 (.D(data_buffer_reg_959__N_3020[896]), .SP(clk_c_enable_1414), 
            .CK(clk_c), .Q(data_buffer_reg[896])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i896.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i897 (.D(data_buffer_reg_959__N_3020[897]), .SP(clk_c_enable_1414), 
            .CK(clk_c), .Q(data_buffer_reg[897])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i897.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i898 (.D(data_buffer_reg_959__N_3020[898]), .SP(clk_c_enable_1414), 
            .CK(clk_c), .Q(data_buffer_reg[898])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i898.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i899 (.D(data_buffer_reg_959__N_3020[899]), .SP(clk_c_enable_1414), 
            .CK(clk_c), .Q(data_buffer_reg[899])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i899.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i900 (.D(data_buffer_reg_959__N_3020[900]), .SP(clk_c_enable_1414), 
            .CK(clk_c), .Q(data_buffer_reg[900])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i900.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i904 (.D(data_buffer_reg_959__N_3020[904]), .SP(clk_c_enable_1414), 
            .CK(clk_c), .Q(data_buffer_reg[904])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i904.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i905 (.D(data_buffer_reg_959__N_3020[905]), .SP(clk_c_enable_1414), 
            .CK(clk_c), .Q(data_buffer_reg[905])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i905.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i906 (.D(data_buffer_reg_959__N_3020[906]), .SP(clk_c_enable_1414), 
            .CK(clk_c), .Q(data_buffer_reg[906])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i906.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i907 (.D(data_buffer_reg_959__N_3020[907]), .SP(clk_c_enable_1414), 
            .CK(clk_c), .Q(data_buffer_reg[907])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i907.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i908 (.D(data_buffer_reg_959__N_3020[908]), .SP(clk_c_enable_1414), 
            .CK(clk_c), .Q(data_buffer_reg[908])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i908.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i912 (.D(data_buffer_reg_959__N_3020[912]), .SP(clk_c_enable_1414), 
            .CK(clk_c), .Q(data_buffer_reg[912])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i912.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i913 (.D(data_buffer_reg_959__N_3020[913]), .SP(clk_c_enable_1414), 
            .CK(clk_c), .Q(data_buffer_reg[913])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i913.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i914 (.D(data_buffer_reg_959__N_3020[914]), .SP(clk_c_enable_1414), 
            .CK(clk_c), .Q(data_buffer_reg[914])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i914.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i915 (.D(data_buffer_reg_959__N_3020[915]), .SP(clk_c_enable_1414), 
            .CK(clk_c), .Q(data_buffer_reg[915])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i915.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i916 (.D(data_buffer_reg_959__N_3020[916]), .SP(clk_c_enable_1414), 
            .CK(clk_c), .Q(data_buffer_reg[916])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i916.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i920 (.D(data_buffer_reg_959__N_3020[920]), .SP(clk_c_enable_1414), 
            .CK(clk_c), .Q(data_buffer_reg[920])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i920.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i921 (.D(data_buffer_reg_959__N_3020[921]), .SP(clk_c_enable_1414), 
            .CK(clk_c), .Q(data_buffer_reg[921])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i921.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i922 (.D(data_buffer_reg_959__N_3020[922]), .SP(clk_c_enable_1414), 
            .CK(clk_c), .Q(data_buffer_reg[922])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i922.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i923 (.D(data_buffer_reg_959__N_3020[923]), .SP(clk_c_enable_1414), 
            .CK(clk_c), .Q(data_buffer_reg[923])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i923.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i924 (.D(data_buffer_reg_959__N_3020[924]), .SP(clk_c_enable_1414), 
            .CK(clk_c), .Q(data_buffer_reg[924])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i924.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i928 (.D(data_buffer_reg_959__N_3020[928]), .SP(clk_c_enable_1414), 
            .CK(clk_c), .Q(data_buffer_reg[928])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i928.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i929 (.D(data_buffer_reg_959__N_3020[929]), .SP(clk_c_enable_1414), 
            .CK(clk_c), .Q(data_buffer_reg[929])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i929.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i930 (.D(data_buffer_reg_959__N_3020[930]), .SP(clk_c_enable_1414), 
            .CK(clk_c), .Q(data_buffer_reg[930])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i930.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i931 (.D(data_buffer_reg_959__N_3020[931]), .SP(clk_c_enable_1414), 
            .CK(clk_c), .Q(data_buffer_reg[931])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i931.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i932 (.D(data_buffer_reg_959__N_3020[932]), .SP(clk_c_enable_1414), 
            .CK(clk_c), .Q(data_buffer_reg[932])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i932.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i936 (.D(data_buffer_reg_959__N_3020[936]), .SP(clk_c_enable_1414), 
            .CK(clk_c), .Q(data_buffer_reg[936])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i936.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i937 (.D(data_buffer_reg_959__N_3020[937]), .SP(clk_c_enable_1414), 
            .CK(clk_c), .Q(data_buffer_reg[937])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i937.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i938 (.D(data_buffer_reg_959__N_3020[938]), .SP(clk_c_enable_1414), 
            .CK(clk_c), .Q(data_buffer_reg[938])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i938.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i939 (.D(data_buffer_reg_959__N_3020[939]), .SP(clk_c_enable_1414), 
            .CK(clk_c), .Q(data_buffer_reg[939])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i939.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i940 (.D(data_buffer_reg_959__N_3020[940]), .SP(clk_c_enable_1414), 
            .CK(clk_c), .Q(data_buffer_reg[940])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i940.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i944 (.D(data_buffer_reg_959__N_3020[944]), .SP(clk_c_enable_1414), 
            .CK(clk_c), .Q(data_buffer_reg[944])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i944.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i945 (.D(data_buffer_reg_959__N_3020[945]), .SP(clk_c_enable_1414), 
            .CK(clk_c), .Q(data_buffer_reg[945])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i945.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i946 (.D(data_buffer_reg_959__N_3020[946]), .SP(clk_c_enable_1414), 
            .CK(clk_c), .Q(data_buffer_reg[946])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i946.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i947 (.D(data_buffer_reg_959__N_3020[947]), .SP(clk_c_enable_1414), 
            .CK(clk_c), .Q(data_buffer_reg[947])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i947.GSR = "ENABLED";
    FD1P3AX data_buffer_reg_i948 (.D(data_buffer_reg_959__N_3020[948]), .SP(clk_c_enable_1414), 
            .CK(clk_c), .Q(data_buffer_reg[948])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i948.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_3_lut_4_lut_rep_494 (.A(data_length_reg[0]), .B(n15), 
         .C(n26793), .D(n25588), .Z(clk_c_enable_1250)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i1_2_lut_3_lut_3_lut_4_lut_rep_494.init = 16'hfef0;
    LUT4 data_buffer_reg_959__I_0_i171_3_lut (.A(data_buffer_reg[178]), .B(\data_buffer[170] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[170])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i171_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i172_3_lut (.A(data_buffer_reg[179]), .B(\data_buffer[171] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[171])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i172_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i1_3_lut (.A(data_buffer_reg[8]), .B(\data_buffer[0] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i1_3_lut.init = 16'hcaca;
    LUT4 i8_4_lut (.A(n15_adj_5036), .B(data_length_reg_c[9]), .C(n14), 
         .D(data_length_reg_c[5]), .Z(n15)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i8_4_lut.init = 16'hfffe;
    LUT4 i6_4_lut (.A(data_length_reg_c[6]), .B(data_length_reg_c[1]), .C(data_length_reg_c[4]), 
         .D(data_length_reg_c[7]), .Z(n15_adj_5036)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i6_4_lut.init = 16'hfffe;
    LUT4 i5_3_lut (.A(data_length_reg_c[3]), .B(data_length_reg_c[2]), .C(data_length_reg_c[8]), 
         .Z(n14)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i5_3_lut.init = 16'hfefe;
    LUT4 i21450_4_lut (.A(cnt[5]), .B(n23729), .C(n21027), .D(cnt[20]), 
         .Z(n24165)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(28[34:52])
    defparam i21450_4_lut.init = 16'h0800;
    LUT4 i20856_4_lut (.A(cnt[4]), .B(cnt[3]), .C(cnt[7]), .D(cnt[6]), 
         .Z(n23723)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i20856_4_lut.init = 16'h8000;
    LUT4 i20933_4_lut (.A(cnt[16]), .B(cnt[2]), .C(cnt[19]), .D(cnt[1]), 
         .Z(n23809)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i20933_4_lut.init = 16'h8000;
    LUT4 i20861_4_lut (.A(cnt[18]), .B(cnt[11]), .C(cnt[0]), .D(cnt[21]), 
         .Z(n23729)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i20861_4_lut.init = 16'h8000;
    LUT4 i9_4_lut (.A(n17), .B(cnt[15]), .C(n16), .D(cnt[10]), .Z(n21027)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(28[34:52])
    defparam i9_4_lut.init = 16'hfffe;
    LUT4 i7_4_lut (.A(cnt[12]), .B(cnt[14]), .C(cnt[23]), .D(cnt[9]), 
         .Z(n17)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(28[34:52])
    defparam i7_4_lut.init = 16'hfffe;
    LUT4 data_buffer_reg_959__I_0_i388_3_lut (.A(data_buffer_reg[395]), .B(\data_buffer[387] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[387])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i388_3_lut.init = 16'hcaca;
    LUT4 i6_4_lut_adj_72 (.A(cnt[8]), .B(cnt[22]), .C(cnt[17]), .D(cnt[13]), 
         .Z(n16)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(28[34:52])
    defparam i6_4_lut_adj_72.init = 16'hfffe;
    LUT4 data_buffer_reg_959__I_0_i173_3_lut (.A(data_buffer_reg[180]), .B(\data_buffer[172] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[172])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i173_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i177_3_lut (.A(data_buffer_reg[184]), .B(\data_buffer[176] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[176])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i177_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i178_3_lut (.A(data_buffer_reg[185]), .B(\data_buffer[177] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[177])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i178_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_341 (.A(data_length_reg[0]), .B(n15), .Z(n25623)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_341.init = 16'heeee;
    LUT4 i9276_2_lut_3_lut_3_lut_4_lut (.A(data_length_reg[0]), .B(n15), 
         .C(n26793), .D(n25588), .Z(n12089)) /* synthesis lut_function=(!(A (C+!(D))+!A ((C+!(D))+!B))) */ ;
    defparam i9276_2_lut_3_lut_3_lut_4_lut.init = 16'h0e00;
    LUT4 i613_2_lut_3_lut (.A(data_length_reg[0]), .B(n15), .C(n3057), 
         .Z(n2025)) /* synthesis lut_function=(A (C)+!A ((C)+!B)) */ ;
    defparam i613_2_lut_3_lut.init = 16'hf1f1;
    LUT4 i1_2_lut_3_lut_3_lut_4_lut (.A(data_length_reg[0]), .B(n15), .C(n26793), 
         .D(n25588), .Z(clk_c_enable_1414)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i1_2_lut_3_lut_3_lut_4_lut.init = 16'hfef0;
    FD1S3IX cnt_1981__i1 (.D(n101[1]), .CK(clk_c), .CD(n25588), .Q(cnt[1])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(19[16:26])
    defparam cnt_1981__i1.GSR = "ENABLED";
    FD1S3IX cnt_1981__i2 (.D(n101[2]), .CK(clk_c), .CD(n25588), .Q(cnt[2])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(19[16:26])
    defparam cnt_1981__i2.GSR = "ENABLED";
    FD1S3IX cnt_1981__i3 (.D(n101[3]), .CK(clk_c), .CD(n25588), .Q(cnt[3])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(19[16:26])
    defparam cnt_1981__i3.GSR = "ENABLED";
    FD1S3IX cnt_1981__i4 (.D(n101[4]), .CK(clk_c), .CD(n25588), .Q(cnt[4])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(19[16:26])
    defparam cnt_1981__i4.GSR = "ENABLED";
    FD1S3IX cnt_1981__i5 (.D(n101[5]), .CK(clk_c), .CD(n25588), .Q(cnt[5])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(19[16:26])
    defparam cnt_1981__i5.GSR = "ENABLED";
    FD1S3IX cnt_1981__i6 (.D(n101[6]), .CK(clk_c), .CD(n25588), .Q(cnt[6])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(19[16:26])
    defparam cnt_1981__i6.GSR = "ENABLED";
    FD1S3IX cnt_1981__i7 (.D(n101[7]), .CK(clk_c), .CD(n25588), .Q(cnt[7])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(19[16:26])
    defparam cnt_1981__i7.GSR = "ENABLED";
    FD1S3IX cnt_1981__i8 (.D(n101[8]), .CK(clk_c), .CD(n25588), .Q(cnt[8])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(19[16:26])
    defparam cnt_1981__i8.GSR = "ENABLED";
    FD1S3IX cnt_1981__i9 (.D(n101[9]), .CK(clk_c), .CD(n25588), .Q(cnt[9])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(19[16:26])
    defparam cnt_1981__i9.GSR = "ENABLED";
    FD1S3IX cnt_1981__i10 (.D(n101[10]), .CK(clk_c), .CD(n25588), .Q(cnt[10])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(19[16:26])
    defparam cnt_1981__i10.GSR = "ENABLED";
    FD1S3IX cnt_1981__i11 (.D(n101[11]), .CK(clk_c), .CD(n25588), .Q(cnt[11])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(19[16:26])
    defparam cnt_1981__i11.GSR = "ENABLED";
    FD1S3IX cnt_1981__i12 (.D(n101[12]), .CK(clk_c), .CD(n25588), .Q(cnt[12])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(19[16:26])
    defparam cnt_1981__i12.GSR = "ENABLED";
    FD1S3IX cnt_1981__i13 (.D(n101[13]), .CK(clk_c), .CD(n25588), .Q(cnt[13])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(19[16:26])
    defparam cnt_1981__i13.GSR = "ENABLED";
    FD1S3IX cnt_1981__i14 (.D(n101[14]), .CK(clk_c), .CD(n25588), .Q(cnt[14])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(19[16:26])
    defparam cnt_1981__i14.GSR = "ENABLED";
    FD1S3IX cnt_1981__i15 (.D(n101[15]), .CK(clk_c), .CD(n25588), .Q(cnt[15])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(19[16:26])
    defparam cnt_1981__i15.GSR = "ENABLED";
    FD1S3IX cnt_1981__i16 (.D(n101[16]), .CK(clk_c), .CD(n25588), .Q(cnt[16])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(19[16:26])
    defparam cnt_1981__i16.GSR = "ENABLED";
    FD1S3IX cnt_1981__i17 (.D(n101[17]), .CK(clk_c), .CD(n25588), .Q(cnt[17])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(19[16:26])
    defparam cnt_1981__i17.GSR = "ENABLED";
    FD1S3IX cnt_1981__i18 (.D(n101[18]), .CK(clk_c), .CD(n25588), .Q(cnt[18])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(19[16:26])
    defparam cnt_1981__i18.GSR = "ENABLED";
    FD1S3IX cnt_1981__i19 (.D(n101[19]), .CK(clk_c), .CD(n25588), .Q(cnt[19])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(19[16:26])
    defparam cnt_1981__i19.GSR = "ENABLED";
    FD1S3IX cnt_1981__i20 (.D(n101[20]), .CK(clk_c), .CD(n25588), .Q(cnt[20])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(19[16:26])
    defparam cnt_1981__i20.GSR = "ENABLED";
    FD1S3IX cnt_1981__i21 (.D(n101[21]), .CK(clk_c), .CD(n25588), .Q(cnt[21])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(19[16:26])
    defparam cnt_1981__i21.GSR = "ENABLED";
    FD1S3IX cnt_1981__i22 (.D(n101[22]), .CK(clk_c), .CD(n25588), .Q(cnt[22])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(19[16:26])
    defparam cnt_1981__i22.GSR = "ENABLED";
    FD1S3IX cnt_1981__i23 (.D(n101[23]), .CK(clk_c), .CD(n25588), .Q(cnt[23])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(19[16:26])
    defparam cnt_1981__i23.GSR = "ENABLED";
    FD1S3AX data_length_reg_1982__i1 (.D(n45[1]), .CK(clk_c), .Q(data_length_reg_c[1])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(29[28:50])
    defparam data_length_reg_1982__i1.GSR = "ENABLED";
    FD1S3AX data_length_reg_1982__i2 (.D(n45[2]), .CK(clk_c), .Q(data_length_reg_c[2])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(29[28:50])
    defparam data_length_reg_1982__i2.GSR = "ENABLED";
    FD1S3AX data_length_reg_1982__i3 (.D(n45[3]), .CK(clk_c), .Q(data_length_reg_c[3])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(29[28:50])
    defparam data_length_reg_1982__i3.GSR = "ENABLED";
    FD1S3AX data_length_reg_1982__i4 (.D(n45[4]), .CK(clk_c), .Q(data_length_reg_c[4])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(29[28:50])
    defparam data_length_reg_1982__i4.GSR = "ENABLED";
    FD1S3AX data_length_reg_1982__i5 (.D(n45[5]), .CK(clk_c), .Q(data_length_reg_c[5])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(29[28:50])
    defparam data_length_reg_1982__i5.GSR = "ENABLED";
    FD1S3AX data_length_reg_1982__i6 (.D(n45[6]), .CK(clk_c), .Q(data_length_reg_c[6])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(29[28:50])
    defparam data_length_reg_1982__i6.GSR = "ENABLED";
    FD1S3AX data_length_reg_1982__i7 (.D(n45[7]), .CK(clk_c), .Q(data_length_reg_c[7])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(29[28:50])
    defparam data_length_reg_1982__i7.GSR = "ENABLED";
    FD1S3AX data_length_reg_1982__i8 (.D(n45[8]), .CK(clk_c), .Q(data_length_reg_c[8])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(29[28:50])
    defparam data_length_reg_1982__i8.GSR = "ENABLED";
    FD1S3AX data_length_reg_1982__i9 (.D(n45[9]), .CK(clk_c), .Q(data_length_reg_c[9])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(29[28:50])
    defparam data_length_reg_1982__i9.GSR = "ENABLED";
    LUT4 data_buffer_reg_959__I_0_i179_3_lut (.A(data_buffer_reg[186]), .B(\data_buffer[178] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[178])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i179_3_lut.init = 16'hcaca;
    FD1P3IX data_buffer_reg_i956 (.D(\data_buffer[956] ), .SP(clk_c_enable_1414), 
            .CD(n12089), .CK(clk_c), .Q(data_buffer_reg[956])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i956.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_3_lut_4_lut_rep_490 (.A(data_length_reg[0]), .B(n15), 
         .C(n26793), .D(n25588), .Z(clk_c_enable_1050)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i1_2_lut_3_lut_3_lut_4_lut_rep_490.init = 16'hfef0;
    LUT4 data_buffer_reg_959__I_0_i180_3_lut (.A(data_buffer_reg[187]), .B(\data_buffer[179] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[179])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i180_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_3_lut_4_lut_rep_492 (.A(data_length_reg[0]), .B(n15), 
         .C(n26793), .D(n25588), .Z(clk_c_enable_1150)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i1_2_lut_3_lut_3_lut_4_lut_rep_492.init = 16'hfef0;
    LUT4 data_buffer_reg_959__I_0_i2_3_lut (.A(data_buffer_reg[9]), .B(\data_buffer[1] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i2_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i3_3_lut (.A(data_buffer_reg[10]), .B(\data_buffer[2] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i3_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i4_3_lut (.A(data_buffer_reg[11]), .B(\data_buffer[3] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i4_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i5_3_lut (.A(data_buffer_reg[12]), .B(\data_buffer[4] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i5_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i9_3_lut (.A(data_buffer_reg[16]), .B(\data_buffer[8] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i9_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i10_3_lut (.A(data_buffer_reg[17]), .B(\data_buffer[9] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i10_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i11_3_lut (.A(data_buffer_reg[18]), .B(\data_buffer[10] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i11_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i12_3_lut (.A(data_buffer_reg[19]), .B(\data_buffer[11] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i12_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i13_3_lut (.A(data_buffer_reg[20]), .B(\data_buffer[12] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i13_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i17_3_lut (.A(data_buffer_reg[24]), .B(\data_buffer[16] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i17_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i18_3_lut (.A(data_buffer_reg[25]), .B(\data_buffer[17] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i18_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i19_3_lut (.A(data_buffer_reg[26]), .B(\data_buffer[18] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i19_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i20_3_lut (.A(data_buffer_reg[27]), .B(\data_buffer[19] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i20_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i21_3_lut (.A(data_buffer_reg[28]), .B(\data_buffer[20] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i21_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i25_3_lut (.A(data_buffer_reg[32]), .B(\data_buffer[24] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i25_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i26_3_lut (.A(data_buffer_reg[33]), .B(\data_buffer[25] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i26_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i27_3_lut (.A(data_buffer_reg[34]), .B(\data_buffer[26] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i27_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i28_3_lut (.A(data_buffer_reg[35]), .B(\data_buffer[27] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i28_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i29_3_lut (.A(data_buffer_reg[36]), .B(\data_buffer[28] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i29_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i33_3_lut (.A(data_buffer_reg[40]), .B(\data_buffer[32] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[32])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i33_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i34_3_lut (.A(data_buffer_reg[41]), .B(\data_buffer[33] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[33])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i34_3_lut.init = 16'hcaca;
    FD1P3IX data_buffer_reg_i955 (.D(\data_buffer[955] ), .SP(clk_c_enable_1414), 
            .CD(n12089), .CK(clk_c), .Q(data_buffer_reg[955])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i955.GSR = "ENABLED";
    LUT4 data_buffer_reg_959__I_0_i35_3_lut (.A(data_buffer_reg[42]), .B(\data_buffer[34] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[34])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i35_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i36_3_lut (.A(data_buffer_reg[43]), .B(\data_buffer[35] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[35])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i36_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i37_3_lut (.A(data_buffer_reg[44]), .B(\data_buffer[36] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[36])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i37_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i41_3_lut (.A(data_buffer_reg[48]), .B(\data_buffer[40] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[40])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i41_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i42_3_lut (.A(data_buffer_reg[49]), .B(\data_buffer[41] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[41])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i42_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i43_3_lut (.A(data_buffer_reg[50]), .B(\data_buffer[42] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[42])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i43_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i44_3_lut (.A(data_buffer_reg[51]), .B(\data_buffer[43] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[43])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i44_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i45_3_lut (.A(data_buffer_reg[52]), .B(\data_buffer[44] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[44])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i45_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i49_3_lut (.A(data_buffer_reg[56]), .B(\data_buffer[48] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[48])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i49_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i50_3_lut (.A(data_buffer_reg[57]), .B(\data_buffer[49] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[49])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i50_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i51_3_lut (.A(data_buffer_reg[58]), .B(\data_buffer[50] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[50])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i51_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i52_3_lut (.A(data_buffer_reg[59]), .B(\data_buffer[51] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[51])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i52_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i53_3_lut (.A(data_buffer_reg[60]), .B(\data_buffer[52] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[52])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i53_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i57_3_lut (.A(data_buffer_reg[64]), .B(\data_buffer[56] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[56])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i57_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i58_3_lut (.A(data_buffer_reg[65]), .B(\data_buffer[57] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[57])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i58_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i59_3_lut (.A(data_buffer_reg[66]), .B(\data_buffer[58] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[58])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i59_3_lut.init = 16'hcaca;
    FD1P3IX data_buffer_reg_i954 (.D(\data_buffer[954] ), .SP(clk_c_enable_1414), 
            .CD(n12089), .CK(clk_c), .Q(data_buffer_reg[954])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i954.GSR = "ENABLED";
    LUT4 data_buffer_reg_959__I_0_i60_3_lut (.A(data_buffer_reg[67]), .B(\data_buffer[59] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[59])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i60_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i61_3_lut (.A(data_buffer_reg[68]), .B(\data_buffer[60] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[60])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i61_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i389_3_lut (.A(data_buffer_reg[396]), .B(\data_buffer[388] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[388])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i389_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i65_3_lut (.A(data_buffer_reg[72]), .B(\data_buffer[64] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[64])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i65_3_lut.init = 16'hcaca;
    FD1P3IX data_buffer_reg_i953 (.D(\data_buffer[953] ), .SP(clk_c_enable_1414), 
            .CD(n12089), .CK(clk_c), .Q(data_buffer_reg[953])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i953.GSR = "ENABLED";
    FD1P3IX data_buffer_reg_i952 (.D(\data_buffer[952] ), .SP(clk_c_enable_1414), 
            .CD(n12089), .CK(clk_c), .Q(data_buffer_reg[952])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=104, LSE_RLINE=113 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(35[10] 39[8])
    defparam data_buffer_reg_i952.GSR = "ENABLED";
    LUT4 data_buffer_reg_959__I_0_i66_3_lut (.A(data_buffer_reg[73]), .B(\data_buffer[65] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[65])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i66_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i181_3_lut (.A(data_buffer_reg[188]), .B(\data_buffer[180] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[180])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i181_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i67_3_lut (.A(data_buffer_reg[74]), .B(\data_buffer[66] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[66])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i67_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i68_3_lut (.A(data_buffer_reg[75]), .B(\data_buffer[67] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[67])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i68_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i69_3_lut (.A(data_buffer_reg[76]), .B(\data_buffer[68] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[68])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i69_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i73_3_lut (.A(data_buffer_reg[80]), .B(\data_buffer[72] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[72])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i73_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i74_3_lut (.A(data_buffer_reg[81]), .B(\data_buffer[73] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[73])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i74_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i75_3_lut (.A(data_buffer_reg[82]), .B(\data_buffer[74] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[74])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i75_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i76_3_lut (.A(data_buffer_reg[83]), .B(\data_buffer[75] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[75])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i76_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i77_3_lut (.A(data_buffer_reg[84]), .B(\data_buffer[76] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[76])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i77_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i81_3_lut (.A(data_buffer_reg[88]), .B(\data_buffer[80] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[80])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i81_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i82_3_lut (.A(data_buffer_reg[89]), .B(\data_buffer[81] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[81])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i82_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i83_3_lut (.A(data_buffer_reg[90]), .B(\data_buffer[82] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[82])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i83_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i84_3_lut (.A(data_buffer_reg[91]), .B(\data_buffer[83] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[83])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i84_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i85_3_lut (.A(data_buffer_reg[92]), .B(\data_buffer[84] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[84])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i85_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i89_3_lut (.A(data_buffer_reg[96]), .B(\data_buffer[88] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[88])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i89_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i185_3_lut (.A(data_buffer_reg[192]), .B(\data_buffer[184] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[184])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i185_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i90_3_lut (.A(data_buffer_reg[97]), .B(\data_buffer[89] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[89])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i90_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i91_3_lut (.A(data_buffer_reg[98]), .B(\data_buffer[90] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[90])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i91_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i186_3_lut (.A(data_buffer_reg[193]), .B(\data_buffer[185] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[185])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i186_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i92_3_lut (.A(data_buffer_reg[99]), .B(\data_buffer[91] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[91])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i92_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i93_3_lut (.A(data_buffer_reg[100]), .B(\data_buffer[92] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[92])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i93_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i97_3_lut (.A(data_buffer_reg[104]), .B(\data_buffer[96] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[96])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i97_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i98_3_lut (.A(data_buffer_reg[105]), .B(\data_buffer[97] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[97])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i98_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i99_3_lut (.A(data_buffer_reg[106]), .B(\data_buffer[98] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[98])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i99_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i100_3_lut (.A(data_buffer_reg[107]), .B(\data_buffer[99] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[99])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i100_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i101_3_lut (.A(data_buffer_reg[108]), .B(\data_buffer[100] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[100])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i101_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i187_3_lut (.A(data_buffer_reg[194]), .B(\data_buffer[186] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[186])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i187_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i105_3_lut (.A(data_buffer_reg[112]), .B(\data_buffer[104] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[104])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i105_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i106_3_lut (.A(data_buffer_reg[113]), .B(\data_buffer[105] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[105])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i106_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i107_3_lut (.A(data_buffer_reg[114]), .B(\data_buffer[106] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[106])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i107_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i108_3_lut (.A(data_buffer_reg[115]), .B(\data_buffer[107] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[107])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i108_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i109_3_lut (.A(data_buffer_reg[116]), .B(\data_buffer[108] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[108])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i109_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i113_3_lut (.A(data_buffer_reg[120]), .B(\data_buffer[112] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[112])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i113_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i114_3_lut (.A(data_buffer_reg[121]), .B(\data_buffer[113] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[113])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i114_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i115_3_lut (.A(data_buffer_reg[122]), .B(\data_buffer[114] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[114])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i115_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i116_3_lut (.A(data_buffer_reg[123]), .B(\data_buffer[115] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[115])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i116_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i117_3_lut (.A(data_buffer_reg[124]), .B(\data_buffer[116] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[116])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i117_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i121_3_lut (.A(data_buffer_reg[128]), .B(\data_buffer[120] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[120])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i121_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i122_3_lut (.A(data_buffer_reg[129]), .B(\data_buffer[121] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[121])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i122_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i123_3_lut (.A(data_buffer_reg[130]), .B(\data_buffer[122] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[122])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i123_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i124_3_lut (.A(data_buffer_reg[131]), .B(\data_buffer[123] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[123])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i124_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i125_3_lut (.A(data_buffer_reg[132]), .B(\data_buffer[124] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[124])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i125_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i129_3_lut (.A(data_buffer_reg[136]), .B(\data_buffer[128] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[128])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i129_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i130_3_lut (.A(data_buffer_reg[137]), .B(\data_buffer[129] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[129])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i130_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i188_3_lut (.A(data_buffer_reg[195]), .B(\data_buffer[187] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[187])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i188_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i131_3_lut (.A(data_buffer_reg[138]), .B(\data_buffer[130] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[130])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i131_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i132_3_lut (.A(data_buffer_reg[139]), .B(\data_buffer[131] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[131])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i132_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i133_3_lut (.A(data_buffer_reg[140]), .B(\data_buffer[132] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[132])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i133_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i137_3_lut (.A(data_buffer_reg[144]), .B(\data_buffer[136] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[136])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i137_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i138_3_lut (.A(data_buffer_reg[145]), .B(\data_buffer[137] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[137])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i138_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_3_lut_4_lut_rep_491 (.A(data_length_reg[0]), .B(n15), 
         .C(n26793), .D(n25588), .Z(clk_c_enable_1100)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i1_2_lut_3_lut_3_lut_4_lut_rep_491.init = 16'hfef0;
    LUT4 data_buffer_reg_959__I_0_i139_3_lut (.A(data_buffer_reg[146]), .B(\data_buffer[138] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[138])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i139_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i140_3_lut (.A(data_buffer_reg[147]), .B(\data_buffer[139] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[139])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i140_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i141_3_lut (.A(data_buffer_reg[148]), .B(\data_buffer[140] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[140])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i141_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i145_3_lut (.A(data_buffer_reg[152]), .B(\data_buffer[144] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[144])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i145_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i146_3_lut (.A(data_buffer_reg[153]), .B(\data_buffer[145] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[145])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i146_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i147_3_lut (.A(data_buffer_reg[154]), .B(\data_buffer[146] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[146])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i147_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i148_3_lut (.A(data_buffer_reg[155]), .B(\data_buffer[147] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[147])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i148_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i149_3_lut (.A(data_buffer_reg[156]), .B(\data_buffer[148] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[148])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i149_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i153_3_lut (.A(data_buffer_reg[160]), .B(\data_buffer[152] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[152])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i153_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i154_3_lut (.A(data_buffer_reg[161]), .B(\data_buffer[153] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[153])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i154_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i155_3_lut (.A(data_buffer_reg[162]), .B(\data_buffer[154] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[154])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i155_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i156_3_lut (.A(data_buffer_reg[163]), .B(\data_buffer[155] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[155])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i156_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i157_3_lut (.A(data_buffer_reg[164]), .B(\data_buffer[156] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[156])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i157_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i189_3_lut (.A(data_buffer_reg[196]), .B(\data_buffer[188] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[188])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i189_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i393_3_lut (.A(data_buffer_reg[400]), .B(\data_buffer[392] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[392])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i393_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i394_3_lut (.A(data_buffer_reg[401]), .B(\data_buffer[393] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[393])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i394_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_3_lut_4_lut_rep_495 (.A(data_length_reg[0]), .B(n15), 
         .C(n26793), .D(n25588), .Z(clk_c_enable_1304)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i1_2_lut_3_lut_3_lut_4_lut_rep_495.init = 16'hfef0;
    LUT4 data_buffer_reg_959__I_0_i395_3_lut (.A(data_buffer_reg[402]), .B(\data_buffer[394] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[394])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i395_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i193_3_lut (.A(data_buffer_reg[200]), .B(\data_buffer[192] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[192])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i193_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i194_3_lut (.A(data_buffer_reg[201]), .B(\data_buffer[193] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[193])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i194_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i195_3_lut (.A(data_buffer_reg[202]), .B(\data_buffer[194] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[194])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i195_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i196_3_lut (.A(data_buffer_reg[203]), .B(\data_buffer[195] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[195])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i196_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i197_3_lut (.A(data_buffer_reg[204]), .B(\data_buffer[196] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[196])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i197_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i201_3_lut (.A(data_buffer_reg[208]), .B(\data_buffer[200] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[200])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i201_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i396_3_lut (.A(data_buffer_reg[403]), .B(\data_buffer[395] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[395])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i396_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i397_3_lut (.A(data_buffer_reg[404]), .B(\data_buffer[396] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[396])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i397_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i202_3_lut (.A(data_buffer_reg[209]), .B(\data_buffer[201] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[201])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i202_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i203_3_lut (.A(data_buffer_reg[210]), .B(\data_buffer[202] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[202])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i203_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i204_3_lut (.A(data_buffer_reg[211]), .B(\data_buffer[203] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[203])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i204_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i205_3_lut (.A(data_buffer_reg[212]), .B(\data_buffer[204] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[204])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i205_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i209_3_lut (.A(data_buffer_reg[216]), .B(\data_buffer[208] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[208])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i209_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i418_3_lut (.A(data_buffer_reg[425]), .B(\data_buffer[417] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[417])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i418_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i419_3_lut (.A(data_buffer_reg[426]), .B(\data_buffer[418] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[418])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i419_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i420_3_lut (.A(data_buffer_reg[427]), .B(\data_buffer[419] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[419])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i420_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i421_3_lut (.A(data_buffer_reg[428]), .B(\data_buffer[420] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[420])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i421_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i401_3_lut (.A(data_buffer_reg[408]), .B(\data_buffer[400] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[400])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i401_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i402_3_lut (.A(data_buffer_reg[409]), .B(\data_buffer[401] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[401])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i402_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i210_3_lut (.A(data_buffer_reg[217]), .B(\data_buffer[209] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[209])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i210_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i211_3_lut (.A(data_buffer_reg[218]), .B(\data_buffer[210] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[210])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i211_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i425_3_lut (.A(data_buffer_reg[432]), .B(\data_buffer[424] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[424])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i425_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i212_3_lut (.A(data_buffer_reg[219]), .B(\data_buffer[211] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[211])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i212_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i426_3_lut (.A(data_buffer_reg[433]), .B(\data_buffer[425] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[425])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i426_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i213_3_lut (.A(data_buffer_reg[220]), .B(\data_buffer[212] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[212])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i213_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i427_3_lut (.A(data_buffer_reg[434]), .B(\data_buffer[426] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[426])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i427_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i403_3_lut (.A(data_buffer_reg[410]), .B(\data_buffer[402] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[402])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i403_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i428_3_lut (.A(data_buffer_reg[435]), .B(\data_buffer[427] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[427])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i428_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i429_3_lut (.A(data_buffer_reg[436]), .B(\data_buffer[428] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[428])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i429_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i217_3_lut (.A(data_buffer_reg[224]), .B(\data_buffer[216] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[216])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i217_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i218_3_lut (.A(data_buffer_reg[225]), .B(\data_buffer[217] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[217])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i218_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i219_3_lut (.A(data_buffer_reg[226]), .B(\data_buffer[218] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[218])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i219_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i220_3_lut (.A(data_buffer_reg[227]), .B(\data_buffer[219] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[219])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i220_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i433_3_lut (.A(data_buffer_reg[440]), .B(\data_buffer[432] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[432])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i433_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i434_3_lut (.A(data_buffer_reg[441]), .B(\data_buffer[433] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[433])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i434_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i221_3_lut (.A(data_buffer_reg[228]), .B(\data_buffer[220] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[220])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i221_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i435_3_lut (.A(data_buffer_reg[442]), .B(\data_buffer[434] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[434])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i435_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i436_3_lut (.A(data_buffer_reg[443]), .B(\data_buffer[435] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[435])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i436_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i437_3_lut (.A(data_buffer_reg[444]), .B(\data_buffer[436] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[436])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i437_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i441_3_lut (.A(data_buffer_reg[448]), .B(\data_buffer[440] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[440])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i441_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i225_3_lut (.A(data_buffer_reg[232]), .B(\data_buffer[224] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[224])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i225_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i226_3_lut (.A(data_buffer_reg[233]), .B(\data_buffer[225] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[225])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i226_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i442_3_lut (.A(data_buffer_reg[449]), .B(\data_buffer[441] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[441])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i442_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i404_3_lut (.A(data_buffer_reg[411]), .B(\data_buffer[403] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[403])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i404_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i227_3_lut (.A(data_buffer_reg[234]), .B(\data_buffer[226] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[226])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i227_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i228_3_lut (.A(data_buffer_reg[235]), .B(\data_buffer[227] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[227])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i228_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i229_3_lut (.A(data_buffer_reg[236]), .B(\data_buffer[228] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[228])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i229_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i233_3_lut (.A(data_buffer_reg[240]), .B(\data_buffer[232] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[232])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i233_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i234_3_lut (.A(data_buffer_reg[241]), .B(\data_buffer[233] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[233])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i234_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i235_3_lut (.A(data_buffer_reg[242]), .B(\data_buffer[234] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[234])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i235_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i443_3_lut (.A(data_buffer_reg[450]), .B(\data_buffer[442] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[442])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i443_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i444_3_lut (.A(data_buffer_reg[451]), .B(\data_buffer[443] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[443])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i444_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i405_3_lut (.A(data_buffer_reg[412]), .B(\data_buffer[404] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[404])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i405_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i445_3_lut (.A(data_buffer_reg[452]), .B(\data_buffer[444] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[444])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i445_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i236_3_lut (.A(data_buffer_reg[243]), .B(\data_buffer[235] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[235])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i236_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i237_3_lut (.A(data_buffer_reg[244]), .B(\data_buffer[236] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[236])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i237_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i409_3_lut (.A(data_buffer_reg[416]), .B(\data_buffer[408] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[408])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i409_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i241_3_lut (.A(data_buffer_reg[248]), .B(\data_buffer[240] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[240])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i241_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i410_3_lut (.A(data_buffer_reg[417]), .B(\data_buffer[409] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[409])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i410_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i242_3_lut (.A(data_buffer_reg[249]), .B(\data_buffer[241] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[241])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i242_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i449_3_lut (.A(data_buffer_reg[456]), .B(\data_buffer[448] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[448])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i449_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i243_3_lut (.A(data_buffer_reg[250]), .B(\data_buffer[242] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[242])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i243_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i450_3_lut (.A(data_buffer_reg[457]), .B(\data_buffer[449] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[449])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i450_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i451_3_lut (.A(data_buffer_reg[458]), .B(\data_buffer[450] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[450])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i451_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i244_3_lut (.A(data_buffer_reg[251]), .B(\data_buffer[243] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[243])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i244_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i452_3_lut (.A(data_buffer_reg[459]), .B(\data_buffer[451] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[451])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i452_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i245_3_lut (.A(data_buffer_reg[252]), .B(\data_buffer[244] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[244])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i245_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i249_3_lut (.A(data_buffer_reg[256]), .B(\data_buffer[248] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[248])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i249_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i453_3_lut (.A(data_buffer_reg[460]), .B(\data_buffer[452] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[452])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i453_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i250_3_lut (.A(data_buffer_reg[257]), .B(\data_buffer[249] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[249])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i250_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i251_3_lut (.A(data_buffer_reg[258]), .B(\data_buffer[250] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[250])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i251_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i252_3_lut (.A(data_buffer_reg[259]), .B(\data_buffer[251] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[251])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i252_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i253_3_lut (.A(data_buffer_reg[260]), .B(\data_buffer[252] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[252])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i253_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i257_3_lut (.A(data_buffer_reg[264]), .B(\data_buffer[256] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[256])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i257_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i258_3_lut (.A(data_buffer_reg[265]), .B(\data_buffer[257] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[257])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i258_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i259_3_lut (.A(data_buffer_reg[266]), .B(\data_buffer[258] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[258])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i259_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i260_3_lut (.A(data_buffer_reg[267]), .B(\data_buffer[259] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[259])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i260_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i261_3_lut (.A(data_buffer_reg[268]), .B(\data_buffer[260] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[260])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i261_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i265_3_lut (.A(data_buffer_reg[272]), .B(\data_buffer[264] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[264])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i265_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i266_3_lut (.A(data_buffer_reg[273]), .B(\data_buffer[265] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[265])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i266_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i267_3_lut (.A(data_buffer_reg[274]), .B(\data_buffer[266] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[266])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i267_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_3_lut_4_lut_rep_486 (.A(data_length_reg[0]), .B(n15), 
         .C(n26793), .D(n25588), .Z(clk_c_enable_849)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i1_2_lut_3_lut_3_lut_4_lut_rep_486.init = 16'hfef0;
    LUT4 data_buffer_reg_959__I_0_i268_3_lut (.A(data_buffer_reg[275]), .B(\data_buffer[267] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[267])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i268_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i269_3_lut (.A(data_buffer_reg[276]), .B(\data_buffer[268] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[268])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i269_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i273_3_lut (.A(data_buffer_reg[280]), .B(\data_buffer[272] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[272])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i273_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i457_3_lut (.A(data_buffer_reg[464]), .B(\data_buffer[456] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[456])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i457_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i274_3_lut (.A(data_buffer_reg[281]), .B(\data_buffer[273] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[273])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i274_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i275_3_lut (.A(data_buffer_reg[282]), .B(\data_buffer[274] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[274])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i275_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i458_3_lut (.A(data_buffer_reg[465]), .B(\data_buffer[457] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[457])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i458_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i276_3_lut (.A(data_buffer_reg[283]), .B(\data_buffer[275] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[275])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i276_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i277_3_lut (.A(data_buffer_reg[284]), .B(\data_buffer[276] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[276])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i277_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i459_3_lut (.A(data_buffer_reg[466]), .B(\data_buffer[458] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[458])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i459_3_lut.init = 16'hcaca;
    CCU2D data_length_reg_1982_add_4_11 (.A0(data_length[8]), .B0(n26793), 
          .C0(data_length_reg_c[8]), .D0(GND_net), .A1(data_length[9]), 
          .B1(n26793), .C1(data_length_reg_c[9]), .D1(GND_net), .CIN(n20546), 
          .S0(n45[8]), .S1(n45[9]));   // g:/fpga/mxo2/system/project/beeper_control.v(29[28:50])
    defparam data_length_reg_1982_add_4_11.INIT0 = 16'h4b8b;
    defparam data_length_reg_1982_add_4_11.INIT1 = 16'h4b8b;
    defparam data_length_reg_1982_add_4_11.INJECT1_0 = "NO";
    defparam data_length_reg_1982_add_4_11.INJECT1_1 = "NO";
    LUT4 data_buffer_reg_959__I_0_i281_3_lut (.A(data_buffer_reg[288]), .B(\data_buffer[280] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[280])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i281_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i460_3_lut (.A(data_buffer_reg[467]), .B(\data_buffer[459] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[459])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i460_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i461_3_lut (.A(data_buffer_reg[468]), .B(\data_buffer[460] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[460])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i461_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i282_3_lut (.A(data_buffer_reg[289]), .B(\data_buffer[281] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[281])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i282_3_lut.init = 16'hcaca;
    CCU2D data_length_reg_1982_add_4_9 (.A0(data_length[6]), .B0(n26793), 
          .C0(data_length_reg_c[6]), .D0(GND_net), .A1(data_length[7]), 
          .B1(n26793), .C1(data_length_reg_c[7]), .D1(GND_net), .CIN(n20545), 
          .COUT(n20546), .S0(n45[6]), .S1(n45[7]));   // g:/fpga/mxo2/system/project/beeper_control.v(29[28:50])
    defparam data_length_reg_1982_add_4_9.INIT0 = 16'h4b8b;
    defparam data_length_reg_1982_add_4_9.INIT1 = 16'h4b8b;
    defparam data_length_reg_1982_add_4_9.INJECT1_0 = "NO";
    defparam data_length_reg_1982_add_4_9.INJECT1_1 = "NO";
    LUT4 data_buffer_reg_959__I_0_i283_3_lut (.A(data_buffer_reg[290]), .B(\data_buffer[282] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[282])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i283_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i284_3_lut (.A(data_buffer_reg[291]), .B(\data_buffer[283] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[283])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i284_3_lut.init = 16'hcaca;
    CCU2D data_length_reg_1982_add_4_7 (.A0(data_length[4]), .B0(n26793), 
          .C0(data_length_reg_c[4]), .D0(GND_net), .A1(data_length[5]), 
          .B1(n26793), .C1(data_length_reg_c[5]), .D1(GND_net), .CIN(n20544), 
          .COUT(n20545), .S0(n45[4]), .S1(n45[5]));   // g:/fpga/mxo2/system/project/beeper_control.v(29[28:50])
    defparam data_length_reg_1982_add_4_7.INIT0 = 16'h4b8b;
    defparam data_length_reg_1982_add_4_7.INIT1 = 16'h4b8b;
    defparam data_length_reg_1982_add_4_7.INJECT1_0 = "NO";
    defparam data_length_reg_1982_add_4_7.INJECT1_1 = "NO";
    CCU2D data_length_reg_1982_add_4_5 (.A0(data_length[2]), .B0(n26793), 
          .C0(data_length_reg_c[2]), .D0(GND_net), .A1(data_length[3]), 
          .B1(n26793), .C1(data_length_reg_c[3]), .D1(GND_net), .CIN(n20543), 
          .COUT(n20544), .S0(n45[2]), .S1(n45[3]));   // g:/fpga/mxo2/system/project/beeper_control.v(29[28:50])
    defparam data_length_reg_1982_add_4_5.INIT0 = 16'h4b8b;
    defparam data_length_reg_1982_add_4_5.INIT1 = 16'h4b8b;
    defparam data_length_reg_1982_add_4_5.INJECT1_0 = "NO";
    defparam data_length_reg_1982_add_4_5.INJECT1_1 = "NO";
    LUT4 data_buffer_reg_959__I_0_i285_3_lut (.A(data_buffer_reg[292]), .B(\data_buffer[284] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[284])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i285_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i289_3_lut (.A(data_buffer_reg[296]), .B(\data_buffer[288] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[288])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i289_3_lut.init = 16'hcaca;
    CCU2D data_length_reg_1982_add_4_3 (.A0(data_length_reg[0]), .B0(n26793), 
          .C0(data_length[0]), .D0(n25562), .A1(data_length[1]), .B1(n26793), 
          .C1(data_length_reg_c[1]), .D1(GND_net), .CIN(n20542), .COUT(n20543), 
          .S0(n45[0]), .S1(n45[1]));   // g:/fpga/mxo2/system/project/beeper_control.v(29[28:50])
    defparam data_length_reg_1982_add_4_3.INIT0 = 16'hd1e2;
    defparam data_length_reg_1982_add_4_3.INIT1 = 16'h4b8b;
    defparam data_length_reg_1982_add_4_3.INJECT1_0 = "NO";
    defparam data_length_reg_1982_add_4_3.INJECT1_1 = "NO";
    LUT4 data_buffer_reg_959__I_0_i465_3_lut (.A(data_buffer_reg[472]), .B(\data_buffer[464] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[464])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i465_3_lut.init = 16'hcaca;
    CCU2D data_length_reg_1982_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n26793), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n20542));   // g:/fpga/mxo2/system/project/beeper_control.v(29[28:50])
    defparam data_length_reg_1982_add_4_1.INIT0 = 16'hF000;
    defparam data_length_reg_1982_add_4_1.INIT1 = 16'h0aaa;
    defparam data_length_reg_1982_add_4_1.INJECT1_0 = "NO";
    defparam data_length_reg_1982_add_4_1.INJECT1_1 = "NO";
    LUT4 data_buffer_reg_959__I_0_i290_3_lut (.A(data_buffer_reg[297]), .B(\data_buffer[289] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[289])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i290_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i466_3_lut (.A(data_buffer_reg[473]), .B(\data_buffer[465] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[465])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i466_3_lut.init = 16'hcaca;
    CCU2D cnt_1981_add_4_25 (.A0(cnt[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n20538), .S0(n101[23]));   // g:/fpga/mxo2/system/project/beeper_control.v(19[16:26])
    defparam cnt_1981_add_4_25.INIT0 = 16'hfaaa;
    defparam cnt_1981_add_4_25.INIT1 = 16'h0000;
    defparam cnt_1981_add_4_25.INJECT1_0 = "NO";
    defparam cnt_1981_add_4_25.INJECT1_1 = "NO";
    LUT4 data_buffer_reg_959__I_0_i291_3_lut (.A(data_buffer_reg[298]), .B(\data_buffer[290] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[290])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i291_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i467_3_lut (.A(data_buffer_reg[474]), .B(\data_buffer[466] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[466])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i467_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i292_3_lut (.A(data_buffer_reg[299]), .B(\data_buffer[291] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[291])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i292_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i293_3_lut (.A(data_buffer_reg[300]), .B(\data_buffer[292] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[292])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i293_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i297_3_lut (.A(data_buffer_reg[304]), .B(\data_buffer[296] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[296])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i297_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i468_3_lut (.A(data_buffer_reg[475]), .B(\data_buffer[467] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[467])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i468_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i298_3_lut (.A(data_buffer_reg[305]), .B(\data_buffer[297] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[297])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i298_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i299_3_lut (.A(data_buffer_reg[306]), .B(\data_buffer[298] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[298])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i299_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i469_3_lut (.A(data_buffer_reg[476]), .B(\data_buffer[468] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[468])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i469_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i473_3_lut (.A(data_buffer_reg[480]), .B(\data_buffer[472] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[472])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i473_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i300_3_lut (.A(data_buffer_reg[307]), .B(\data_buffer[299] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[299])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i300_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i301_3_lut (.A(data_buffer_reg[308]), .B(\data_buffer[300] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[300])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i301_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i305_3_lut (.A(data_buffer_reg[312]), .B(\data_buffer[304] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[304])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i305_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i306_3_lut (.A(data_buffer_reg[313]), .B(\data_buffer[305] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[305])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i306_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i307_3_lut (.A(data_buffer_reg[314]), .B(\data_buffer[306] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[306])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i307_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i308_3_lut (.A(data_buffer_reg[315]), .B(\data_buffer[307] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[307])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i308_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i309_3_lut (.A(data_buffer_reg[316]), .B(\data_buffer[308] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[308])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i309_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i313_3_lut (.A(data_buffer_reg[320]), .B(\data_buffer[312] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[312])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i313_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i474_3_lut (.A(data_buffer_reg[481]), .B(\data_buffer[473] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[473])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i474_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i314_3_lut (.A(data_buffer_reg[321]), .B(\data_buffer[313] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[313])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i314_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i315_3_lut (.A(data_buffer_reg[322]), .B(\data_buffer[314] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[314])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i315_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i316_3_lut (.A(data_buffer_reg[323]), .B(\data_buffer[315] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[315])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i316_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i475_3_lut (.A(data_buffer_reg[482]), .B(\data_buffer[474] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[474])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i475_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i317_3_lut (.A(data_buffer_reg[324]), .B(\data_buffer[316] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[316])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i317_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i476_3_lut (.A(data_buffer_reg[483]), .B(\data_buffer[475] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[475])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i476_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i321_3_lut (.A(data_buffer_reg[328]), .B(\data_buffer[320] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[320])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i321_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i322_3_lut (.A(data_buffer_reg[329]), .B(\data_buffer[321] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[321])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i322_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i477_3_lut (.A(data_buffer_reg[484]), .B(\data_buffer[476] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[476])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i477_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i481_3_lut (.A(data_buffer_reg[488]), .B(\data_buffer[480] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[480])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i481_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i323_3_lut (.A(data_buffer_reg[330]), .B(\data_buffer[322] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[322])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i323_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i324_3_lut (.A(data_buffer_reg[331]), .B(\data_buffer[323] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[323])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i324_3_lut.init = 16'hcaca;
    CCU2D cnt_1981_add_4_23 (.A0(cnt[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[22]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n20537), .COUT(n20538), .S0(n101[21]), .S1(n101[22]));   // g:/fpga/mxo2/system/project/beeper_control.v(19[16:26])
    defparam cnt_1981_add_4_23.INIT0 = 16'hfaaa;
    defparam cnt_1981_add_4_23.INIT1 = 16'hfaaa;
    defparam cnt_1981_add_4_23.INJECT1_0 = "NO";
    defparam cnt_1981_add_4_23.INJECT1_1 = "NO";
    LUT4 data_buffer_reg_959__I_0_i325_3_lut (.A(data_buffer_reg[332]), .B(\data_buffer[324] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[324])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i325_3_lut.init = 16'hcaca;
    CCU2D cnt_1981_add_4_21 (.A0(cnt[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[20]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n20536), .COUT(n20537), .S0(n101[19]), .S1(n101[20]));   // g:/fpga/mxo2/system/project/beeper_control.v(19[16:26])
    defparam cnt_1981_add_4_21.INIT0 = 16'hfaaa;
    defparam cnt_1981_add_4_21.INIT1 = 16'hfaaa;
    defparam cnt_1981_add_4_21.INJECT1_0 = "NO";
    defparam cnt_1981_add_4_21.INJECT1_1 = "NO";
    LUT4 data_buffer_reg_959__I_0_i482_3_lut (.A(data_buffer_reg[489]), .B(\data_buffer[481] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[481])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i482_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i329_3_lut (.A(data_buffer_reg[336]), .B(\data_buffer[328] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[328])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i329_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i330_3_lut (.A(data_buffer_reg[337]), .B(\data_buffer[329] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[329])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i330_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i331_3_lut (.A(data_buffer_reg[338]), .B(\data_buffer[330] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[330])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i331_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i332_3_lut (.A(data_buffer_reg[339]), .B(\data_buffer[331] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[331])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i332_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i483_3_lut (.A(data_buffer_reg[490]), .B(\data_buffer[482] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[482])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i483_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i484_3_lut (.A(data_buffer_reg[491]), .B(\data_buffer[483] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[483])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i484_3_lut.init = 16'hcaca;
    CCU2D cnt_1981_add_4_19 (.A0(cnt[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n20535), .COUT(n20536), .S0(n101[17]), .S1(n101[18]));   // g:/fpga/mxo2/system/project/beeper_control.v(19[16:26])
    defparam cnt_1981_add_4_19.INIT0 = 16'hfaaa;
    defparam cnt_1981_add_4_19.INIT1 = 16'hfaaa;
    defparam cnt_1981_add_4_19.INJECT1_0 = "NO";
    defparam cnt_1981_add_4_19.INJECT1_1 = "NO";
    LUT4 data_buffer_reg_959__I_0_i485_3_lut (.A(data_buffer_reg[492]), .B(\data_buffer[484] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[484])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i485_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i333_3_lut (.A(data_buffer_reg[340]), .B(\data_buffer[332] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[332])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i333_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i489_3_lut (.A(data_buffer_reg[496]), .B(\data_buffer[488] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[488])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i489_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i337_3_lut (.A(data_buffer_reg[344]), .B(\data_buffer[336] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[336])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i337_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i338_3_lut (.A(data_buffer_reg[345]), .B(\data_buffer[337] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[337])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i338_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i490_3_lut (.A(data_buffer_reg[497]), .B(\data_buffer[489] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[489])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i490_3_lut.init = 16'hcaca;
    CCU2D cnt_1981_add_4_17 (.A0(cnt[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n20534), .COUT(n20535), .S0(n101[15]), .S1(n101[16]));   // g:/fpga/mxo2/system/project/beeper_control.v(19[16:26])
    defparam cnt_1981_add_4_17.INIT0 = 16'hfaaa;
    defparam cnt_1981_add_4_17.INIT1 = 16'hfaaa;
    defparam cnt_1981_add_4_17.INJECT1_0 = "NO";
    defparam cnt_1981_add_4_17.INJECT1_1 = "NO";
    CCU2D cnt_1981_add_4_15 (.A0(cnt[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n20533), .COUT(n20534), .S0(n101[13]), .S1(n101[14]));   // g:/fpga/mxo2/system/project/beeper_control.v(19[16:26])
    defparam cnt_1981_add_4_15.INIT0 = 16'hfaaa;
    defparam cnt_1981_add_4_15.INIT1 = 16'hfaaa;
    defparam cnt_1981_add_4_15.INJECT1_0 = "NO";
    defparam cnt_1981_add_4_15.INJECT1_1 = "NO";
    LUT4 data_buffer_reg_959__I_0_i339_3_lut (.A(data_buffer_reg[346]), .B(\data_buffer[338] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[338])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i339_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i491_3_lut (.A(data_buffer_reg[498]), .B(\data_buffer[490] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[490])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i491_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i340_3_lut (.A(data_buffer_reg[347]), .B(\data_buffer[339] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[339])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i340_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i492_3_lut (.A(data_buffer_reg[499]), .B(\data_buffer[491] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[491])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i492_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i341_3_lut (.A(data_buffer_reg[348]), .B(\data_buffer[340] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[340])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i341_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i345_3_lut (.A(data_buffer_reg[352]), .B(\data_buffer[344] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[344])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i345_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i493_3_lut (.A(data_buffer_reg[500]), .B(\data_buffer[492] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[492])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i493_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i346_3_lut (.A(data_buffer_reg[353]), .B(\data_buffer[345] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[345])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i346_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i497_3_lut (.A(data_buffer_reg[504]), .B(\data_buffer[496] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[496])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i497_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i498_3_lut (.A(data_buffer_reg[505]), .B(\data_buffer[497] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[497])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i498_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i347_3_lut (.A(data_buffer_reg[354]), .B(\data_buffer[346] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[346])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i347_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i348_3_lut (.A(data_buffer_reg[355]), .B(\data_buffer[347] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[347])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i348_3_lut.init = 16'hcaca;
    CCU2D cnt_1981_add_4_13 (.A0(cnt[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n20532), .COUT(n20533), .S0(n101[11]), .S1(n101[12]));   // g:/fpga/mxo2/system/project/beeper_control.v(19[16:26])
    defparam cnt_1981_add_4_13.INIT0 = 16'hfaaa;
    defparam cnt_1981_add_4_13.INIT1 = 16'hfaaa;
    defparam cnt_1981_add_4_13.INJECT1_0 = "NO";
    defparam cnt_1981_add_4_13.INJECT1_1 = "NO";
    CCU2D cnt_1981_add_4_11 (.A0(cnt[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n20531), .COUT(n20532), .S0(n101[9]), .S1(n101[10]));   // g:/fpga/mxo2/system/project/beeper_control.v(19[16:26])
    defparam cnt_1981_add_4_11.INIT0 = 16'hfaaa;
    defparam cnt_1981_add_4_11.INIT1 = 16'hfaaa;
    defparam cnt_1981_add_4_11.INJECT1_0 = "NO";
    defparam cnt_1981_add_4_11.INJECT1_1 = "NO";
    LUT4 data_buffer_reg_959__I_0_i499_3_lut (.A(data_buffer_reg[506]), .B(\data_buffer[498] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[498])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i499_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i500_3_lut (.A(data_buffer_reg[507]), .B(\data_buffer[499] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[499])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i500_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i501_3_lut (.A(data_buffer_reg[508]), .B(\data_buffer[500] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[500])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i501_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i349_3_lut (.A(data_buffer_reg[356]), .B(\data_buffer[348] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[348])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i349_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i353_3_lut (.A(data_buffer_reg[360]), .B(\data_buffer[352] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[352])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i353_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i354_3_lut (.A(data_buffer_reg[361]), .B(\data_buffer[353] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[353])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i354_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i355_3_lut (.A(data_buffer_reg[362]), .B(\data_buffer[354] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[354])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i355_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i356_3_lut (.A(data_buffer_reg[363]), .B(\data_buffer[355] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[355])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i356_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i357_3_lut (.A(data_buffer_reg[364]), .B(\data_buffer[356] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[356])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i357_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i505_3_lut (.A(data_buffer_reg[512]), .B(\data_buffer[504] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[504])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i505_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i361_3_lut (.A(data_buffer_reg[368]), .B(\data_buffer[360] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[360])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i361_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i362_3_lut (.A(data_buffer_reg[369]), .B(\data_buffer[361] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[361])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i362_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i506_3_lut (.A(data_buffer_reg[513]), .B(\data_buffer[505] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[505])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i506_3_lut.init = 16'hcaca;
    CCU2D cnt_1981_add_4_9 (.A0(cnt[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n20530), 
          .COUT(n20531), .S0(n101[7]), .S1(n101[8]));   // g:/fpga/mxo2/system/project/beeper_control.v(19[16:26])
    defparam cnt_1981_add_4_9.INIT0 = 16'hfaaa;
    defparam cnt_1981_add_4_9.INIT1 = 16'hfaaa;
    defparam cnt_1981_add_4_9.INJECT1_0 = "NO";
    defparam cnt_1981_add_4_9.INJECT1_1 = "NO";
    CCU2D cnt_1981_add_4_7 (.A0(cnt[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n20529), 
          .COUT(n20530), .S0(n101[5]), .S1(n101[6]));   // g:/fpga/mxo2/system/project/beeper_control.v(19[16:26])
    defparam cnt_1981_add_4_7.INIT0 = 16'hfaaa;
    defparam cnt_1981_add_4_7.INIT1 = 16'hfaaa;
    defparam cnt_1981_add_4_7.INJECT1_0 = "NO";
    defparam cnt_1981_add_4_7.INJECT1_1 = "NO";
    CCU2D cnt_1981_add_4_5 (.A0(cnt[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n20528), 
          .COUT(n20529), .S0(n101[3]), .S1(n101[4]));   // g:/fpga/mxo2/system/project/beeper_control.v(19[16:26])
    defparam cnt_1981_add_4_5.INIT0 = 16'hfaaa;
    defparam cnt_1981_add_4_5.INIT1 = 16'hfaaa;
    defparam cnt_1981_add_4_5.INJECT1_0 = "NO";
    defparam cnt_1981_add_4_5.INJECT1_1 = "NO";
    LUT4 data_buffer_reg_959__I_0_i507_3_lut (.A(data_buffer_reg[514]), .B(\data_buffer[506] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[506])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i507_3_lut.init = 16'hcaca;
    CCU2D cnt_1981_add_4_3 (.A0(cnt[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n20527), 
          .COUT(n20528), .S0(n101[1]), .S1(n101[2]));   // g:/fpga/mxo2/system/project/beeper_control.v(19[16:26])
    defparam cnt_1981_add_4_3.INIT0 = 16'hfaaa;
    defparam cnt_1981_add_4_3.INIT1 = 16'hfaaa;
    defparam cnt_1981_add_4_3.INJECT1_0 = "NO";
    defparam cnt_1981_add_4_3.INJECT1_1 = "NO";
    LUT4 data_buffer_reg_959__I_0_i363_3_lut (.A(data_buffer_reg[370]), .B(\data_buffer[362] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[362])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i363_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i508_3_lut (.A(data_buffer_reg[515]), .B(\data_buffer[507] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[507])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i508_3_lut.init = 16'hcaca;
    CCU2D cnt_1981_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n20527), .S1(n101[0]));   // g:/fpga/mxo2/system/project/beeper_control.v(19[16:26])
    defparam cnt_1981_add_4_1.INIT0 = 16'hF000;
    defparam cnt_1981_add_4_1.INIT1 = 16'h0555;
    defparam cnt_1981_add_4_1.INJECT1_0 = "NO";
    defparam cnt_1981_add_4_1.INJECT1_1 = "NO";
    LUT4 data_buffer_reg_959__I_0_i364_3_lut (.A(data_buffer_reg[371]), .B(\data_buffer[363] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[363])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i364_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i509_3_lut (.A(data_buffer_reg[516]), .B(\data_buffer[508] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[508])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i509_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i365_3_lut (.A(data_buffer_reg[372]), .B(\data_buffer[364] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[364])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i365_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i369_3_lut (.A(data_buffer_reg[376]), .B(\data_buffer[368] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[368])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i369_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i370_3_lut (.A(data_buffer_reg[377]), .B(\data_buffer[369] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[369])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i370_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i513_3_lut (.A(data_buffer_reg[520]), .B(\data_buffer[512] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[512])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i513_3_lut.init = 16'hcaca;
    LUT4 i21451_3_lut_rep_306 (.A(n24165), .B(n23723), .C(n23809), .Z(n25588)) /* synthesis lut_function=(A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(28[34:52])
    defparam i21451_3_lut_rep_306.init = 16'h8080;
    LUT4 data_buffer_reg_959__I_0_i514_3_lut (.A(data_buffer_reg[521]), .B(\data_buffer[513] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[513])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i514_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i515_3_lut (.A(data_buffer_reg[522]), .B(\data_buffer[514] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[514])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i515_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i516_3_lut (.A(data_buffer_reg[523]), .B(\data_buffer[515] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[515])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i516_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i371_3_lut (.A(data_buffer_reg[378]), .B(\data_buffer[370] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[370])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i371_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i517_3_lut (.A(data_buffer_reg[524]), .B(\data_buffer[516] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[516])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i517_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i521_3_lut (.A(data_buffer_reg[528]), .B(\data_buffer[520] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[520])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i521_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i372_3_lut (.A(data_buffer_reg[379]), .B(\data_buffer[371] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[371])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i372_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i522_3_lut (.A(data_buffer_reg[529]), .B(\data_buffer[521] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[521])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i522_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i373_3_lut (.A(data_buffer_reg[380]), .B(\data_buffer[372] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[372])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i373_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i523_3_lut (.A(data_buffer_reg[530]), .B(\data_buffer[522] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[522])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i523_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i524_3_lut (.A(data_buffer_reg[531]), .B(\data_buffer[523] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[523])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i524_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i525_3_lut (.A(data_buffer_reg[532]), .B(\data_buffer[524] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[524])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i525_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i377_3_lut (.A(data_buffer_reg[384]), .B(\data_buffer[376] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[376])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i377_3_lut.init = 16'hcaca;
    LUT4 i21436_2_lut_rep_280_2_lut_4_lut (.A(n24165), .B(n23723), .C(n23809), 
         .D(n25623), .Z(n25562)) /* synthesis lut_function=(!(A (B (C (D))))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(28[34:52])
    defparam i21436_2_lut_rep_280_2_lut_4_lut.init = 16'h7fff;
    LUT4 data_buffer_reg_959__I_0_i529_3_lut (.A(data_buffer_reg[536]), .B(\data_buffer[528] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[528])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i529_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i530_3_lut (.A(data_buffer_reg[537]), .B(\data_buffer[529] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[529])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i530_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i531_3_lut (.A(data_buffer_reg[538]), .B(\data_buffer[530] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[530])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i531_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i532_3_lut (.A(data_buffer_reg[539]), .B(\data_buffer[531] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[531])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i532_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i533_3_lut (.A(data_buffer_reg[540]), .B(\data_buffer[532] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[532])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i533_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i537_3_lut (.A(data_buffer_reg[544]), .B(\data_buffer[536] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[536])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i537_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i538_3_lut (.A(data_buffer_reg[545]), .B(\data_buffer[537] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[537])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i538_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i378_3_lut (.A(data_buffer_reg[385]), .B(\data_buffer[377] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[377])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i378_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i379_3_lut (.A(data_buffer_reg[386]), .B(\data_buffer[378] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[378])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i379_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i380_3_lut (.A(data_buffer_reg[387]), .B(\data_buffer[379] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[379])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i380_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i381_3_lut (.A(data_buffer_reg[388]), .B(\data_buffer[380] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[380])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i381_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i411_3_lut (.A(data_buffer_reg[418]), .B(\data_buffer[410] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[410])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i411_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i412_3_lut (.A(data_buffer_reg[419]), .B(\data_buffer[411] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[411])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i412_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i413_3_lut (.A(data_buffer_reg[420]), .B(\data_buffer[412] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[412])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i413_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i385_3_lut (.A(data_buffer_reg[392]), .B(\data_buffer[384] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[384])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i385_3_lut.init = 16'hcaca;
    LUT4 data_buffer_reg_959__I_0_i386_3_lut (.A(data_buffer_reg[393]), .B(\data_buffer[385] ), 
         .C(n26793), .Z(data_buffer_reg_959__N_3020[385])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(37[10] 39[8])
    defparam data_buffer_reg_959__I_0_i386_3_lut.init = 16'hcaca;
    Beeper Beeper_inst (.GND_net(GND_net), .n3057(n3057), .\data_buffer_reg[3] (data_buffer_reg[3]), 
           .\data_buffer_reg[1] (data_buffer_reg[1]), .\data_buffer_reg[2] (data_buffer_reg[2]), 
           .\data_buffer_reg[4] (data_buffer_reg[4]), .piano_out_c(piano_out_c), 
           .clk_c(clk_c), .\data_buffer_reg[0] (data_buffer_reg[0]), .n2025(n2025)) /* synthesis syn_module_defined=1 */ ;   // g:/fpga/mxo2/system/project/beeper_control.v(49[8] 55[2])
    
endmodule
//
// Verilog Description of module Beeper
//

module Beeper (GND_net, n3057, \data_buffer_reg[3] , \data_buffer_reg[1] , 
            \data_buffer_reg[2] , \data_buffer_reg[4] , piano_out_c, clk_c, 
            \data_buffer_reg[0] , n2025) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output n3057;
    input \data_buffer_reg[3] ;
    input \data_buffer_reg[1] ;
    input \data_buffer_reg[2] ;
    input \data_buffer_reg[4] ;
    output piano_out_c;
    input clk_c;
    input \data_buffer_reg[0] ;
    input n2025;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // g:/fpga/mxo2/system/project/system_top.v(2[15:18])
    
    wire n20518;
    wire [17:0]time_cnt;   // g:/fpga/mxo2/system/project/beeper.v(39[12:20])
    wire [17:0]n3038;
    
    wire n25828, n25827, n15, n30;
    wire [15:0]time_end;   // g:/fpga/mxo2/system/project/beeper.v(10[12:20])
    
    wire n25831, n25830, piano_out_N_5017, n20517, n25837, n25836, 
        n24628, n15_adj_5032, n30_adj_5033, n20516, n25778, n25779, 
        n20515, n7, n5794, n15_adj_5034, n25540;
    wire [17:0]n77;
    
    wire n20514, n25793, n25794, n20513, n24633, n24634, n20512, 
        n20511, n20510, n23797, n36, n23795, n23793, n30_adj_5035, 
        n23533, n23690, n25662, n25541, n24796, n24627, n24795, 
        n20570, n20569, n20568, n20567, n20566, n20565, n20564, 
        n20563, n20562, n25782, n25781, n25813, n25812, n25816, 
        n25815, n25819, n25818;
    
    CCU2D add_1033_19 (.A0(time_cnt[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n20518), .S0(n3038[17]), .S1(n3057));   // g:/fpga/mxo2/system/project/beeper.v(46[14:32])
    defparam add_1033_19.INIT0 = 16'h5555;
    defparam add_1033_19.INIT1 = 16'h0000;
    defparam add_1033_19.INJECT1_0 = "NO";
    defparam add_1033_19.INJECT1_1 = "NO";
    LUT4 tone_4__I_0_26_Mux_2_i31_then_4_lut (.A(\data_buffer_reg[3] ), .B(\data_buffer_reg[1] ), 
         .C(\data_buffer_reg[2] ), .D(\data_buffer_reg[4] ), .Z(n25828)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C (D))+!B ((D)+!C))) */ ;
    defparam tone_4__I_0_26_Mux_2_i31_then_4_lut.init = 16'hfb8b;
    LUT4 tone_4__I_0_26_Mux_2_i31_else_4_lut (.A(\data_buffer_reg[3] ), .B(\data_buffer_reg[1] ), 
         .C(\data_buffer_reg[2] ), .D(\data_buffer_reg[4] ), .Z(n25827)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C+(D)))+!A (B ((D)+!C)+!B !(D))) */ ;
    defparam tone_4__I_0_26_Mux_2_i31_else_4_lut.init = 16'hee3d;
    PFUMX tone_4__I_0_26_Mux_8_i31 (.BLUT(n15), .ALUT(n30), .C0(\data_buffer_reg[4] ), 
          .Z(time_end[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=49, LSE_RLINE=55 */ ;
    LUT4 tone_4__I_0_26_Mux_9_i31_then_4_lut (.A(\data_buffer_reg[1] ), .B(\data_buffer_reg[2] ), 
         .C(\data_buffer_reg[4] ), .D(\data_buffer_reg[3] ), .Z(n25831)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(D))) */ ;
    defparam tone_4__I_0_26_Mux_9_i31_then_4_lut.init = 16'hfdee;
    LUT4 tone_4__I_0_26_Mux_9_i31_else_4_lut (.A(\data_buffer_reg[1] ), .B(\data_buffer_reg[2] ), 
         .C(\data_buffer_reg[4] ), .D(\data_buffer_reg[3] ), .Z(n25830)) /* synthesis lut_function=(A (B (C+(D))+!B ((D)+!C))+!A (B (C (D)+!C !(D))+!B (C+!(D)))) */ ;
    defparam tone_4__I_0_26_Mux_9_i31_else_4_lut.init = 16'hfa97;
    FD1S3AX piano_out_23 (.D(piano_out_N_5017), .CK(clk_c), .Q(piano_out_c)) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=49, LSE_RLINE=55 */ ;   // g:/fpga/mxo2/system/project/beeper.v(57[11] 61[5])
    defparam piano_out_23.GSR = "ENABLED";
    CCU2D add_1033_17 (.A0(time_cnt[15]), .B0(time_end[15]), .C0(GND_net), 
          .D0(GND_net), .A1(time_cnt[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n20517), .COUT(n20518), .S0(n3038[15]), 
          .S1(n3038[16]));   // g:/fpga/mxo2/system/project/beeper.v(46[14:32])
    defparam add_1033_17.INIT0 = 16'h5999;
    defparam add_1033_17.INIT1 = 16'h5555;
    defparam add_1033_17.INJECT1_0 = "NO";
    defparam add_1033_17.INJECT1_1 = "NO";
    LUT4 tone_4__I_0_26_Mux_12_i31_then_4_lut (.A(\data_buffer_reg[4] ), .B(\data_buffer_reg[1] ), 
         .C(\data_buffer_reg[2] ), .D(\data_buffer_reg[3] ), .Z(n25837)) /* synthesis lut_function=(A (B (C+(D))+!B ((D)+!C))+!A (B (C (D))+!B (C+!(D)))) */ ;
    defparam tone_4__I_0_26_Mux_12_i31_then_4_lut.init = 16'hfa93;
    LUT4 tone_4__I_0_26_Mux_12_i31_else_4_lut (.A(\data_buffer_reg[4] ), .B(\data_buffer_reg[1] ), 
         .C(\data_buffer_reg[2] ), .D(\data_buffer_reg[3] ), .Z(n25836)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)+!C !(D)))) */ ;
    defparam tone_4__I_0_26_Mux_12_i31_else_4_lut.init = 16'hfacb;
    LUT4 n1_bdd_4_lut_21634 (.A(\data_buffer_reg[0] ), .B(\data_buffer_reg[2] ), 
         .C(\data_buffer_reg[4] ), .D(\data_buffer_reg[1] ), .Z(n24628)) /* synthesis lut_function=(A (B+(C (D)+!C !(D)))+!A (B (C)+!B !(C))) */ ;
    defparam n1_bdd_4_lut_21634.init = 16'he9cb;
    PFUMX tone_4__I_0_26_Mux_1_i31 (.BLUT(n15_adj_5032), .ALUT(n30_adj_5033), 
          .C0(\data_buffer_reg[4] ), .Z(time_end[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=49, LSE_RLINE=55 */ ;
    CCU2D add_1033_15 (.A0(time_cnt[13]), .B0(time_end[13]), .C0(GND_net), 
          .D0(GND_net), .A1(time_cnt[14]), .B1(time_end[14]), .C1(GND_net), 
          .D1(GND_net), .CIN(n20516), .COUT(n20517), .S0(n3038[13]), 
          .S1(n3038[14]));   // g:/fpga/mxo2/system/project/beeper.v(46[14:32])
    defparam add_1033_15.INIT0 = 16'h5999;
    defparam add_1033_15.INIT1 = 16'h5999;
    defparam add_1033_15.INJECT1_0 = "NO";
    defparam add_1033_15.INJECT1_1 = "NO";
    PFUMX i22159 (.BLUT(n25778), .ALUT(n25779), .C0(\data_buffer_reg[0] ), 
          .Z(time_end[14]));
    CCU2D add_1033_13 (.A0(time_cnt[11]), .B0(time_end[11]), .C0(GND_net), 
          .D0(GND_net), .A1(time_cnt[12]), .B1(time_end[12]), .C1(GND_net), 
          .D1(GND_net), .CIN(n20515), .COUT(n20516), .S0(n3038[11]), 
          .S1(n3038[12]));   // g:/fpga/mxo2/system/project/beeper.v(46[14:32])
    defparam add_1033_13.INIT0 = 16'h5999;
    defparam add_1033_13.INIT1 = 16'h5999;
    defparam add_1033_13.INJECT1_0 = "NO";
    defparam add_1033_13.INJECT1_1 = "NO";
    PFUMX tone_4__I_0_26_Mux_6_i15 (.BLUT(n7), .ALUT(n5794), .C0(\data_buffer_reg[3] ), 
          .Z(n15_adj_5034)) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=8, LSE_RCOL=2, LSE_LLINE=49, LSE_RLINE=55 */ ;
    LUT4 n3_bdd_4_lut_22142 (.A(\data_buffer_reg[0] ), .B(\data_buffer_reg[4] ), 
         .C(\data_buffer_reg[3] ), .D(\data_buffer_reg[1] ), .Z(n25540)) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)))+!A (B (C+(D))+!B ((D)+!C))) */ ;
    defparam n3_bdd_4_lut_22142.init = 16'hdfe3;
    FD1S3IX time_cnt_1987__i0 (.D(n77[0]), .CK(clk_c), .CD(n2025), .Q(time_cnt[0])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/beeper.v(49[15:30])
    defparam time_cnt_1987__i0.GSR = "ENABLED";
    CCU2D add_1033_11 (.A0(time_cnt[9]), .B0(time_end[9]), .C0(GND_net), 
          .D0(GND_net), .A1(time_cnt[10]), .B1(time_end[10]), .C1(GND_net), 
          .D1(GND_net), .CIN(n20514), .COUT(n20515), .S0(n3038[9]), 
          .S1(n3038[10]));   // g:/fpga/mxo2/system/project/beeper.v(46[14:32])
    defparam add_1033_11.INIT0 = 16'h5999;
    defparam add_1033_11.INIT1 = 16'h5999;
    defparam add_1033_11.INJECT1_0 = "NO";
    defparam add_1033_11.INJECT1_1 = "NO";
    PFUMX i22169 (.BLUT(n25793), .ALUT(n25794), .C0(\data_buffer_reg[3] ), 
          .Z(time_end[10]));
    CCU2D add_1033_9 (.A0(time_cnt[7]), .B0(time_end[7]), .C0(GND_net), 
          .D0(GND_net), .A1(time_cnt[8]), .B1(time_end[8]), .C1(GND_net), 
          .D1(GND_net), .CIN(n20513), .COUT(n20514), .S0(n3038[7]), 
          .S1(n3038[8]));   // g:/fpga/mxo2/system/project/beeper.v(46[14:32])
    defparam add_1033_9.INIT0 = 16'h5999;
    defparam add_1033_9.INIT1 = 16'h5999;
    defparam add_1033_9.INJECT1_0 = "NO";
    defparam add_1033_9.INJECT1_1 = "NO";
    LUT4 data_buffer_reg_3__bdd_4_lut (.A(\data_buffer_reg[3] ), .B(\data_buffer_reg[2] ), 
         .C(\data_buffer_reg[4] ), .D(\data_buffer_reg[0] ), .Z(n24633)) /* synthesis lut_function=(A ((C+!(D))+!B)+!A (B (C)+!B (C+!(D)))) */ ;
    defparam data_buffer_reg_3__bdd_4_lut.init = 16'hf2fb;
    LUT4 data_buffer_reg_3__bdd_3_lut_21637 (.A(\data_buffer_reg[3] ), .B(\data_buffer_reg[2] ), 
         .C(\data_buffer_reg[0] ), .Z(n24634)) /* synthesis lut_function=(A+((C)+!B)) */ ;
    defparam data_buffer_reg_3__bdd_3_lut_21637.init = 16'hfbfb;
    CCU2D add_1033_7 (.A0(time_cnt[5]), .B0(time_end[5]), .C0(GND_net), 
          .D0(GND_net), .A1(n15_adj_5034), .B1(\data_buffer_reg[4] ), 
          .C1(time_cnt[6]), .D1(GND_net), .CIN(n20512), .COUT(n20513), 
          .S0(n3038[5]), .S1(n3038[6]));   // g:/fpga/mxo2/system/project/beeper.v(46[14:32])
    defparam add_1033_7.INIT0 = 16'h5999;
    defparam add_1033_7.INIT1 = 16'he1e1;
    defparam add_1033_7.INJECT1_0 = "NO";
    defparam add_1033_7.INJECT1_1 = "NO";
    CCU2D add_1033_5 (.A0(time_cnt[3]), .B0(time_end[3]), .C0(GND_net), 
          .D0(GND_net), .A1(time_cnt[4]), .B1(time_end[4]), .C1(GND_net), 
          .D1(GND_net), .CIN(n20511), .COUT(n20512), .S0(n3038[3]), 
          .S1(n3038[4]));   // g:/fpga/mxo2/system/project/beeper.v(46[14:32])
    defparam add_1033_5.INIT0 = 16'h5999;
    defparam add_1033_5.INIT1 = 16'h5999;
    defparam add_1033_5.INJECT1_0 = "NO";
    defparam add_1033_5.INJECT1_1 = "NO";
    CCU2D add_1033_3 (.A0(time_cnt[1]), .B0(time_end[1]), .C0(GND_net), 
          .D0(GND_net), .A1(time_cnt[2]), .B1(time_end[2]), .C1(GND_net), 
          .D1(GND_net), .CIN(n20510), .COUT(n20511), .S0(n3038[1]), 
          .S1(n3038[2]));   // g:/fpga/mxo2/system/project/beeper.v(46[14:32])
    defparam add_1033_3.INIT0 = 16'h5999;
    defparam add_1033_3.INIT1 = 16'h5999;
    defparam add_1033_3.INJECT1_0 = "NO";
    defparam add_1033_3.INJECT1_1 = "NO";
    CCU2D add_1033_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(time_cnt[0]), .B1(time_end[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n20510), .S1(n3038[0]));   // g:/fpga/mxo2/system/project/beeper.v(46[14:32])
    defparam add_1033_1.INIT0 = 16'h0000;
    defparam add_1033_1.INIT1 = 16'h5999;
    defparam add_1033_1.INJECT1_0 = "NO";
    defparam add_1033_1.INJECT1_1 = "NO";
    LUT4 i21552_4_lut_4_lut_then_4_lut (.A(\data_buffer_reg[0] ), .B(\data_buffer_reg[2] ), 
         .C(\data_buffer_reg[4] ), .D(\data_buffer_reg[1] ), .Z(n25794)) /* synthesis lut_function=(A (B (C+(D))+!B (C+!(D)))+!A (B+(C+!(D)))) */ ;   // g:/fpga/mxo2/system/project/beeper.v(13[2] 36[9])
    defparam i21552_4_lut_4_lut_then_4_lut.init = 16'hfcf7;
    LUT4 i21552_4_lut_4_lut_else_4_lut (.A(\data_buffer_reg[0] ), .B(\data_buffer_reg[2] ), 
         .C(\data_buffer_reg[4] ), .D(\data_buffer_reg[1] ), .Z(n25793)) /* synthesis lut_function=(A (D)+!A (B (C+(D))+!B !(C))) */ ;   // g:/fpga/mxo2/system/project/beeper.v(13[2] 36[9])
    defparam i21552_4_lut_4_lut_else_4_lut.init = 16'hef41;
    FD1S3IX time_cnt_1987__i1 (.D(n77[1]), .CK(clk_c), .CD(n2025), .Q(time_cnt[1])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/beeper.v(49[15:30])
    defparam time_cnt_1987__i1.GSR = "ENABLED";
    FD1S3IX time_cnt_1987__i2 (.D(n77[2]), .CK(clk_c), .CD(n2025), .Q(time_cnt[2])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/beeper.v(49[15:30])
    defparam time_cnt_1987__i2.GSR = "ENABLED";
    FD1S3IX time_cnt_1987__i3 (.D(n77[3]), .CK(clk_c), .CD(n2025), .Q(time_cnt[3])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/beeper.v(49[15:30])
    defparam time_cnt_1987__i3.GSR = "ENABLED";
    FD1S3IX time_cnt_1987__i4 (.D(n77[4]), .CK(clk_c), .CD(n2025), .Q(time_cnt[4])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/beeper.v(49[15:30])
    defparam time_cnt_1987__i4.GSR = "ENABLED";
    FD1S3IX time_cnt_1987__i5 (.D(n77[5]), .CK(clk_c), .CD(n2025), .Q(time_cnt[5])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/beeper.v(49[15:30])
    defparam time_cnt_1987__i5.GSR = "ENABLED";
    FD1S3IX time_cnt_1987__i6 (.D(n77[6]), .CK(clk_c), .CD(n2025), .Q(time_cnt[6])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/beeper.v(49[15:30])
    defparam time_cnt_1987__i6.GSR = "ENABLED";
    FD1S3IX time_cnt_1987__i7 (.D(n77[7]), .CK(clk_c), .CD(n2025), .Q(time_cnt[7])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/beeper.v(49[15:30])
    defparam time_cnt_1987__i7.GSR = "ENABLED";
    FD1S3IX time_cnt_1987__i8 (.D(n77[8]), .CK(clk_c), .CD(n2025), .Q(time_cnt[8])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/beeper.v(49[15:30])
    defparam time_cnt_1987__i8.GSR = "ENABLED";
    FD1S3IX time_cnt_1987__i9 (.D(n77[9]), .CK(clk_c), .CD(n2025), .Q(time_cnt[9])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/beeper.v(49[15:30])
    defparam time_cnt_1987__i9.GSR = "ENABLED";
    FD1S3IX time_cnt_1987__i10 (.D(n77[10]), .CK(clk_c), .CD(n2025), .Q(time_cnt[10])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/beeper.v(49[15:30])
    defparam time_cnt_1987__i10.GSR = "ENABLED";
    FD1S3IX time_cnt_1987__i11 (.D(n77[11]), .CK(clk_c), .CD(n2025), .Q(time_cnt[11])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/beeper.v(49[15:30])
    defparam time_cnt_1987__i11.GSR = "ENABLED";
    FD1S3IX time_cnt_1987__i12 (.D(n77[12]), .CK(clk_c), .CD(n2025), .Q(time_cnt[12])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/beeper.v(49[15:30])
    defparam time_cnt_1987__i12.GSR = "ENABLED";
    FD1S3IX time_cnt_1987__i13 (.D(n77[13]), .CK(clk_c), .CD(n2025), .Q(time_cnt[13])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/beeper.v(49[15:30])
    defparam time_cnt_1987__i13.GSR = "ENABLED";
    FD1S3IX time_cnt_1987__i14 (.D(n77[14]), .CK(clk_c), .CD(n2025), .Q(time_cnt[14])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/beeper.v(49[15:30])
    defparam time_cnt_1987__i14.GSR = "ENABLED";
    FD1S3IX time_cnt_1987__i15 (.D(n77[15]), .CK(clk_c), .CD(n2025), .Q(time_cnt[15])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/beeper.v(49[15:30])
    defparam time_cnt_1987__i15.GSR = "ENABLED";
    FD1S3IX time_cnt_1987__i16 (.D(n77[16]), .CK(clk_c), .CD(n2025), .Q(time_cnt[16])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/beeper.v(49[15:30])
    defparam time_cnt_1987__i16.GSR = "ENABLED";
    FD1S3IX time_cnt_1987__i17 (.D(n77[17]), .CK(clk_c), .CD(n2025), .Q(time_cnt[17])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/beeper.v(49[15:30])
    defparam time_cnt_1987__i17.GSR = "ENABLED";
    LUT4 piano_out_I_0_4_lut (.A(piano_out_c), .B(n23797), .C(n36), .D(n23795), 
         .Z(piano_out_N_5017)) /* synthesis lut_function=(A (B+((D)+!C))+!A !(B+((D)+!C))) */ ;   // g:/fpga/mxo2/system/project/beeper.v(59[11] 61[5])
    defparam piano_out_I_0_4_lut.init = 16'haa9a;
    LUT4 i20921_4_lut (.A(n3038[8]), .B(n3038[3]), .C(n3038[4]), .D(n3038[17]), 
         .Z(n23797)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20921_4_lut.init = 16'hfffe;
    LUT4 i17_4_lut (.A(n23793), .B(n3038[12]), .C(n30_adj_5035), .D(n23533), 
         .Z(n36)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i17_4_lut.init = 16'h0010;
    LUT4 i20919_4_lut (.A(n3038[10]), .B(n3038[0]), .C(n3038[7]), .D(n3038[15]), 
         .Z(n23795)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20919_4_lut.init = 16'hfffe;
    LUT4 i20917_4_lut (.A(n3038[6]), .B(n3038[11]), .C(n3038[16]), .D(n3038[9]), 
         .Z(n23793)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20917_4_lut.init = 16'hfffe;
    LUT4 i11_4_lut (.A(n23690), .B(n3038[13]), .C(\data_buffer_reg[4] ), 
         .D(n25662), .Z(n30_adj_5035)) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i11_4_lut.init = 16'h1110;
    LUT4 i20696_2_lut (.A(n3038[1]), .B(n3038[2]), .Z(n23533)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i20696_2_lut.init = 16'heeee;
    LUT4 i20826_2_lut (.A(n3038[14]), .B(n3038[5]), .Z(n23690)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i20826_2_lut.init = 16'heeee;
    LUT4 n3_bdd_4_lut_4_lut (.A(\data_buffer_reg[1] ), .B(\data_buffer_reg[3] ), 
         .C(\data_buffer_reg[4] ), .D(\data_buffer_reg[0] ), .Z(n25541)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A ((C+(D))+!B)) */ ;   // g:/fpga/mxo2/system/project/beeper.v(13[2] 36[9])
    defparam n3_bdd_4_lut_4_lut.init = 16'hffd1;
    LUT4 i13597_2_lut_3_lut_3_lut (.A(\data_buffer_reg[1] ), .B(\data_buffer_reg[3] ), 
         .C(\data_buffer_reg[2] ), .Z(n30)) /* synthesis lut_function=((B+(C))+!A) */ ;   // g:/fpga/mxo2/system/project/beeper.v(13[2] 36[9])
    defparam i13597_2_lut_3_lut_3_lut.init = 16'hfdfd;
    LUT4 i13325_4_lut_4_lut (.A(\data_buffer_reg[0] ), .B(\data_buffer_reg[2] ), 
         .C(\data_buffer_reg[1] ), .D(\data_buffer_reg[3] ), .Z(n30_adj_5033)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A ((C+(D))+!B)) */ ;   // g:/fpga/mxo2/system/project/beeper.v(13[2] 36[9])
    defparam i13325_4_lut_4_lut.init = 16'hffd1;
    LUT4 data_buffer_reg_4__bdd_4_lut_4_lut (.A(\data_buffer_reg[0] ), .B(\data_buffer_reg[3] ), 
         .C(\data_buffer_reg[2] ), .D(\data_buffer_reg[1] ), .Z(n24796)) /* synthesis lut_function=(A (B (D)+!B !(C (D)+!C !(D)))+!A (B ((D)+!C)+!B !(C (D)))) */ ;   // g:/fpga/mxo2/system/project/beeper.v(13[2] 36[9])
    defparam data_buffer_reg_4__bdd_4_lut_4_lut.init = 16'hcf35;
    LUT4 n1_bdd_4_lut_21625_4_lut_4_lut (.A(\data_buffer_reg[0] ), .B(\data_buffer_reg[2] ), 
         .C(\data_buffer_reg[4] ), .D(\data_buffer_reg[1] ), .Z(n24627)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A (C+!(D))) */ ;   // g:/fpga/mxo2/system/project/beeper.v(13[2] 36[9])
    defparam n1_bdd_4_lut_21625_4_lut_4_lut.init = 16'hf0fd;
    LUT4 data_buffer_reg_4__bdd_3_lut_4_lut (.A(\data_buffer_reg[0] ), .B(\data_buffer_reg[1] ), 
         .C(\data_buffer_reg[3] ), .D(\data_buffer_reg[2] ), .Z(n24795)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;
    defparam data_buffer_reg_4__bdd_3_lut_4_lut.init = 16'hfef0;
    LUT4 i13290_4_lut_4_lut_4_lut_4_lut (.A(\data_buffer_reg[0] ), .B(\data_buffer_reg[1] ), 
         .C(\data_buffer_reg[2] ), .D(\data_buffer_reg[3] ), .Z(n15)) /* synthesis lut_function=(!(A (C (D))+!A !(B+(C+!(D))))) */ ;
    defparam i13290_4_lut_4_lut_4_lut_4_lut.init = 16'h5eff;
    LUT4 tone_4__I_0_26_Mux_6_i7_3_lut_3_lut_3_lut (.A(\data_buffer_reg[0] ), 
         .B(\data_buffer_reg[1] ), .C(\data_buffer_reg[2] ), .Z(n7)) /* synthesis lut_function=(A (C)+!A (B+!(C))) */ ;
    defparam tone_4__I_0_26_Mux_6_i7_3_lut_3_lut_3_lut.init = 16'he5e5;
    LUT4 i2999_3_lut_3_lut (.A(\data_buffer_reg[0] ), .B(\data_buffer_reg[1] ), 
         .C(\data_buffer_reg[2] ), .Z(n5794)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B)) */ ;   // g:/fpga/mxo2/system/project/beeper.v(13[2] 36[9])
    defparam i2999_3_lut_3_lut.init = 16'h9393;
    LUT4 tone_4__I_0_26_Mux_14_i31_3_lut_then_4_lut (.A(\data_buffer_reg[4] ), 
         .B(\data_buffer_reg[1] ), .C(\data_buffer_reg[2] ), .D(\data_buffer_reg[3] ), 
         .Z(n25779)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A !(C+(D))) */ ;   // g:/fpga/mxo2/system/project/beeper.v(13[2] 36[9])
    defparam tone_4__I_0_26_Mux_14_i31_3_lut_then_4_lut.init = 16'haa85;
    PFUMX i21628 (.BLUT(n24634), .ALUT(n24633), .C0(\data_buffer_reg[1] ), 
          .Z(time_end[7]));
    LUT4 i1_2_lut_rep_380_3_lut_4_lut (.A(\data_buffer_reg[3] ), .B(\data_buffer_reg[1] ), 
         .C(\data_buffer_reg[0] ), .D(\data_buffer_reg[2] ), .Z(n25662)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_380_3_lut_4_lut.init = 16'hfffe;
    CCU2D time_cnt_1987_add_4_19 (.A0(time_cnt[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n20570), .S0(n77[17]));   // g:/fpga/mxo2/system/project/beeper.v(49[15:30])
    defparam time_cnt_1987_add_4_19.INIT0 = 16'hfaaa;
    defparam time_cnt_1987_add_4_19.INIT1 = 16'h0000;
    defparam time_cnt_1987_add_4_19.INJECT1_0 = "NO";
    defparam time_cnt_1987_add_4_19.INJECT1_1 = "NO";
    CCU2D time_cnt_1987_add_4_17 (.A0(time_cnt[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(time_cnt[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n20569), .COUT(n20570), .S0(n77[15]), .S1(n77[16]));   // g:/fpga/mxo2/system/project/beeper.v(49[15:30])
    defparam time_cnt_1987_add_4_17.INIT0 = 16'hfaaa;
    defparam time_cnt_1987_add_4_17.INIT1 = 16'hfaaa;
    defparam time_cnt_1987_add_4_17.INJECT1_0 = "NO";
    defparam time_cnt_1987_add_4_17.INJECT1_1 = "NO";
    CCU2D time_cnt_1987_add_4_15 (.A0(time_cnt[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(time_cnt[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n20568), .COUT(n20569), .S0(n77[13]), .S1(n77[14]));   // g:/fpga/mxo2/system/project/beeper.v(49[15:30])
    defparam time_cnt_1987_add_4_15.INIT0 = 16'hfaaa;
    defparam time_cnt_1987_add_4_15.INIT1 = 16'hfaaa;
    defparam time_cnt_1987_add_4_15.INJECT1_0 = "NO";
    defparam time_cnt_1987_add_4_15.INJECT1_1 = "NO";
    CCU2D time_cnt_1987_add_4_13 (.A0(time_cnt[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(time_cnt[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n20567), .COUT(n20568), .S0(n77[11]), .S1(n77[12]));   // g:/fpga/mxo2/system/project/beeper.v(49[15:30])
    defparam time_cnt_1987_add_4_13.INIT0 = 16'hfaaa;
    defparam time_cnt_1987_add_4_13.INIT1 = 16'hfaaa;
    defparam time_cnt_1987_add_4_13.INJECT1_0 = "NO";
    defparam time_cnt_1987_add_4_13.INJECT1_1 = "NO";
    LUT4 tone_4__I_0_26_Mux_14_i31_3_lut_else_4_lut (.A(\data_buffer_reg[4] ), 
         .B(\data_buffer_reg[1] ), .C(\data_buffer_reg[2] ), .D(\data_buffer_reg[3] ), 
         .Z(n25778)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A !(B (C+(D))+!B (D))) */ ;   // g:/fpga/mxo2/system/project/beeper.v(13[2] 36[9])
    defparam tone_4__I_0_26_Mux_14_i31_3_lut_else_4_lut.init = 16'haa95;
    CCU2D time_cnt_1987_add_4_11 (.A0(time_cnt[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(time_cnt[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n20566), .COUT(n20567), .S0(n77[9]), .S1(n77[10]));   // g:/fpga/mxo2/system/project/beeper.v(49[15:30])
    defparam time_cnt_1987_add_4_11.INIT0 = 16'hfaaa;
    defparam time_cnt_1987_add_4_11.INIT1 = 16'hfaaa;
    defparam time_cnt_1987_add_4_11.INJECT1_0 = "NO";
    defparam time_cnt_1987_add_4_11.INJECT1_1 = "NO";
    CCU2D time_cnt_1987_add_4_9 (.A0(time_cnt[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(time_cnt[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n20565), .COUT(n20566), .S0(n77[7]), .S1(n77[8]));   // g:/fpga/mxo2/system/project/beeper.v(49[15:30])
    defparam time_cnt_1987_add_4_9.INIT0 = 16'hfaaa;
    defparam time_cnt_1987_add_4_9.INIT1 = 16'hfaaa;
    defparam time_cnt_1987_add_4_9.INJECT1_0 = "NO";
    defparam time_cnt_1987_add_4_9.INJECT1_1 = "NO";
    CCU2D time_cnt_1987_add_4_7 (.A0(time_cnt[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(time_cnt[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n20564), .COUT(n20565), .S0(n77[5]), .S1(n77[6]));   // g:/fpga/mxo2/system/project/beeper.v(49[15:30])
    defparam time_cnt_1987_add_4_7.INIT0 = 16'hfaaa;
    defparam time_cnt_1987_add_4_7.INIT1 = 16'hfaaa;
    defparam time_cnt_1987_add_4_7.INJECT1_0 = "NO";
    defparam time_cnt_1987_add_4_7.INJECT1_1 = "NO";
    CCU2D time_cnt_1987_add_4_5 (.A0(time_cnt[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(time_cnt[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n20563), .COUT(n20564), .S0(n77[3]), .S1(n77[4]));   // g:/fpga/mxo2/system/project/beeper.v(49[15:30])
    defparam time_cnt_1987_add_4_5.INIT0 = 16'hfaaa;
    defparam time_cnt_1987_add_4_5.INIT1 = 16'hfaaa;
    defparam time_cnt_1987_add_4_5.INJECT1_0 = "NO";
    defparam time_cnt_1987_add_4_5.INJECT1_1 = "NO";
    PFUMX i21626 (.BLUT(n24628), .ALUT(n24627), .C0(\data_buffer_reg[3] ), 
          .Z(time_end[11]));
    CCU2D time_cnt_1987_add_4_3 (.A0(time_cnt[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(time_cnt[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n20562), .COUT(n20563), .S0(n77[1]), .S1(n77[2]));   // g:/fpga/mxo2/system/project/beeper.v(49[15:30])
    defparam time_cnt_1987_add_4_3.INIT0 = 16'hfaaa;
    defparam time_cnt_1987_add_4_3.INIT1 = 16'hfaaa;
    defparam time_cnt_1987_add_4_3.INJECT1_0 = "NO";
    defparam time_cnt_1987_add_4_3.INJECT1_1 = "NO";
    CCU2D time_cnt_1987_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(time_cnt[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n20562), .S1(n77[0]));   // g:/fpga/mxo2/system/project/beeper.v(49[15:30])
    defparam time_cnt_1987_add_4_1.INIT0 = 16'hF000;
    defparam time_cnt_1987_add_4_1.INIT1 = 16'h0555;
    defparam time_cnt_1987_add_4_1.INJECT1_0 = "NO";
    defparam time_cnt_1987_add_4_1.INJECT1_1 = "NO";
    LUT4 tone_4__I_0_26_Mux_13_i31_3_lut_then_4_lut (.A(\data_buffer_reg[4] ), 
         .B(\data_buffer_reg[1] ), .C(\data_buffer_reg[3] ), .D(\data_buffer_reg[2] ), 
         .Z(n25782)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A !(C (D)+!C !(D))) */ ;   // g:/fpga/mxo2/system/project/beeper.v(13[2] 36[9])
    defparam tone_4__I_0_26_Mux_13_i31_3_lut_then_4_lut.init = 16'hadf0;
    LUT4 tone_4__I_0_26_Mux_13_i31_3_lut_else_4_lut (.A(\data_buffer_reg[4] ), 
         .B(\data_buffer_reg[1] ), .C(\data_buffer_reg[3] ), .D(\data_buffer_reg[2] ), 
         .Z(n25781)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A !(B (C (D)+!C !(D))+!B (D))) */ ;   // g:/fpga/mxo2/system/project/beeper.v(13[2] 36[9])
    defparam tone_4__I_0_26_Mux_13_i31_3_lut_else_4_lut.init = 16'hacf1;
    LUT4 tone_4__I_0_26_Mux_1_i15_4_lut_4_lut_4_lut (.A(\data_buffer_reg[2] ), 
         .B(\data_buffer_reg[0] ), .C(\data_buffer_reg[1] ), .D(\data_buffer_reg[3] ), 
         .Z(n15_adj_5032)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B (C (D))+!B (C+(D))))) */ ;   // g:/fpga/mxo2/system/project/beeper.v(13[2] 36[9])
    defparam tone_4__I_0_26_Mux_1_i15_4_lut_4_lut_4_lut.init = 16'h04e5;
    PFUMX i22143 (.BLUT(n25541), .ALUT(n25540), .C0(\data_buffer_reg[2] ), 
          .Z(time_end[0]));
    PFUMX i22161 (.BLUT(n25781), .ALUT(n25782), .C0(\data_buffer_reg[0] ), 
          .Z(time_end[13]));
    LUT4 n24647_bdd_3_lut_then_4_lut (.A(\data_buffer_reg[3] ), .B(\data_buffer_reg[4] ), 
         .C(\data_buffer_reg[0] ), .D(\data_buffer_reg[2] ), .Z(n25813)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+(D))+!B (C))) */ ;
    defparam n24647_bdd_3_lut_then_4_lut.init = 16'hded8;
    LUT4 n24647_bdd_3_lut_else_4_lut (.A(\data_buffer_reg[3] ), .B(\data_buffer_reg[4] ), 
         .C(\data_buffer_reg[0] ), .D(\data_buffer_reg[2] ), .Z(n25812)) /* synthesis lut_function=(A (B)+!A (B ((D)+!C)+!B !(C (D)))) */ ;
    defparam n24647_bdd_3_lut_else_4_lut.init = 16'hcd9d;
    LUT4 tone_4__I_0_26_Mux_15_i31_3_lut_4_lut_then_1_lut (.A(\data_buffer_reg[4] ), 
         .Z(n25816)) /* synthesis lut_function=(A) */ ;   // g:/fpga/mxo2/system/project/beeper.v(57[37:49])
    defparam tone_4__I_0_26_Mux_15_i31_3_lut_4_lut_then_1_lut.init = 16'haaaa;
    PFUMX i21709 (.BLUT(n24796), .ALUT(n24795), .C0(\data_buffer_reg[4] ), 
          .Z(time_end[3]));
    LUT4 tone_4__I_0_26_Mux_15_i31_3_lut_4_lut_else_1_lut (.A(\data_buffer_reg[0] ), 
         .B(\data_buffer_reg[2] ), .C(\data_buffer_reg[4] ), .D(\data_buffer_reg[1] ), 
         .Z(n25815)) /* synthesis lut_function=(A (B (C (D)))+!A (B (C (D))+!B !(C+(D)))) */ ;   // g:/fpga/mxo2/system/project/beeper.v(57[37:49])
    defparam tone_4__I_0_26_Mux_15_i31_3_lut_4_lut_else_1_lut.init = 16'hc001;
    PFUMX i22198 (.BLUT(n25836), .ALUT(n25837), .C0(\data_buffer_reg[0] ), 
          .Z(time_end[12]));
    LUT4 n25525_bdd_3_lut_then_4_lut (.A(\data_buffer_reg[3] ), .B(\data_buffer_reg[4] ), 
         .C(\data_buffer_reg[1] ), .D(\data_buffer_reg[2] ), .Z(n25819)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;
    defparam n25525_bdd_3_lut_then_4_lut.init = 16'hfaca;
    LUT4 n25525_bdd_3_lut_else_4_lut (.A(\data_buffer_reg[3] ), .B(\data_buffer_reg[4] ), 
         .C(\data_buffer_reg[1] ), .D(\data_buffer_reg[2] ), .Z(n25818)) /* synthesis lut_function=(A (B+(D))+!A (B (C (D)+!C !(D))+!B !(C+(D)))) */ ;
    defparam n25525_bdd_3_lut_else_4_lut.init = 16'hea8d;
    PFUMX i22194 (.BLUT(n25830), .ALUT(n25831), .C0(\data_buffer_reg[0] ), 
          .Z(time_end[9]));
    PFUMX i22192 (.BLUT(n25827), .ALUT(n25828), .C0(\data_buffer_reg[0] ), 
          .Z(time_end[2]));
    PFUMX i22186 (.BLUT(n25818), .ALUT(n25819), .C0(\data_buffer_reg[0] ), 
          .Z(time_end[5]));
    PFUMX i22184 (.BLUT(n25815), .ALUT(n25816), .C0(\data_buffer_reg[3] ), 
          .Z(time_end[15]));
    PFUMX i22182 (.BLUT(n25812), .ALUT(n25813), .C0(\data_buffer_reg[1] ), 
          .Z(time_end[4]));
    
endmodule
//
// Verilog Description of module uart_top
//

module uart_top (\data_buffer[432] , clk_c, clk_c_enable_659, \data_buffer[424] , 
            \data_buffer[0] , \data_buffer[956] , \data_buffer[948] , 
            \data_buffer[955] , \data_buffer[947] , \data_buffer[954] , 
            \data_buffer[946] , \data_buffer[953] , \data_buffer[945] , 
            \data_buffer[952] , \data_buffer[944] , \data_buffer[940] , 
            \data_buffer[939] , \data_buffer[938] , \data_buffer[937] , 
            \data_buffer[936] , \data_buffer[932] , \data_buffer[931] , 
            \data_buffer[930] , \data_buffer[929] , \data_buffer[928] , 
            \data_buffer[924] , \data_buffer[923] , \data_buffer[922] , 
            \data_buffer[921] , \data_buffer[920] , \data_buffer[916] , 
            \data_buffer[915] , \data_buffer[914] , \data_buffer[913] , 
            \data_buffer[912] , \data_buffer[908] , \data_buffer[907] , 
            \data_buffer[906] , \data_buffer[905] , \data_buffer[904] , 
            \data_buffer[900] , \data_buffer[899] , \data_buffer[898] , 
            \data_buffer[897] , \data_buffer[896] , \data_buffer[892] , 
            \data_buffer[891] , \data_buffer[428] , \data_buffer[420] , 
            \data_buffer[427] , \data_buffer[419] , \data_buffer[890] , 
            \data_buffer[889] , \data_buffer[888] , \data_buffer[884] , 
            \data_buffer[883] , \data_buffer[882] , \data_buffer[881] , 
            \data_buffer[880] , \data_buffer[876] , \data_buffer[875] , 
            \data_buffer[874] , \data_buffer[873] , \data_buffer[872] , 
            \data_buffer[868] , \data_buffer[867] , \data_buffer[866] , 
            \data_buffer[865] , \data_buffer[864] , \data_buffer[860] , 
            \data_buffer[859] , \data_buffer[858] , \data_buffer[857] , 
            \data_buffer[856] , \data_buffer[852] , \data_buffer[851] , 
            \data_buffer[850] , \data_buffer[849] , \data_buffer[848] , 
            \data_buffer[844] , \data_buffer[843] , \data_buffer[842] , 
            \data_buffer[841] , \data_buffer[840] , \data_buffer[836] , 
            \data_buffer[835] , \data_buffer[834] , \data_buffer[833] , 
            \data_buffer[832] , \data_buffer[828] , \data_buffer[827] , 
            \data_buffer[826] , \data_buffer[825] , \data_buffer[824] , 
            \data_buffer[820] , \data_buffer[819] , \data_buffer[818] , 
            \data_buffer[817] , \data_buffer[816] , \data_buffer[812] , 
            \data_buffer[811] , \data_buffer[810] , \data_buffer[809] , 
            \data_buffer[808] , \data_buffer[804] , \data_buffer[803] , 
            \data_buffer[802] , \data_buffer[801] , \data_buffer[800] , 
            \data_buffer[796] , \data_buffer[795] , \data_buffer[794] , 
            \data_buffer[793] , \data_buffer[792] , n26780, \data_buffer[788] , 
            \data_buffer[787] , \data_buffer[786] , \data_buffer[785] , 
            \data_buffer[784] , \data_buffer[780] , \data_buffer[779] , 
            \data_buffer[778] , \data_buffer[777] , \data_buffer[776] , 
            \data_buffer[772] , \data_buffer[771] , \data_buffer[770] , 
            \data_buffer[769] , \data_buffer[768] , \data_buffer[764] , 
            \data_buffer[763] , \data_buffer[762] , \data_buffer[761] , 
            \data_buffer[760] , \data_buffer[756] , \data_buffer[755] , 
            \data_buffer[754] , \data_buffer[753] , \data_buffer[752] , 
            \data_buffer[748] , \data_buffer[747] , \data_buffer[746] , 
            \data_buffer[745] , \data_buffer[744] , \data_buffer[740] , 
            \data_buffer[739] , \data_buffer[738] , \data_buffer[737] , 
            \data_buffer[736] , \data_buffer[732] , \data_buffer[731] , 
            \data_buffer[730] , \data_buffer[729] , \data_buffer[728] , 
            \data_buffer[724] , \data_buffer[723] , \data_buffer[722] , 
            \data_buffer[721] , \data_buffer[720] , \data_buffer[716] , 
            \data_buffer[715] , \data_buffer[714] , \data_buffer[713] , 
            \data_buffer[712] , \data_buffer[708] , \data_buffer[707] , 
            \data_buffer[706] , \data_buffer[705] , \data_buffer[704] , 
            \data_buffer[700] , \data_buffer[699] , \data_buffer[698] , 
            \data_buffer[697] , \data_buffer[696] , \data_buffer[692] , 
            \data_buffer[691] , \data_buffer[690] , \data_buffer[689] , 
            \data_buffer[688] , \data_buffer[684] , \data_buffer[683] , 
            \data_buffer[682] , \data_buffer[681] , \data_buffer[680] , 
            \data_buffer[676] , \data_buffer[675] , \data_buffer[674] , 
            \data_buffer[673] , \data_buffer[672] , \data_buffer[668] , 
            \data_buffer[667] , \data_buffer[666] , \data_buffer[665] , 
            \data_buffer[664] , \data_buffer[660] , \data_buffer[659] , 
            \data_buffer[658] , \data_buffer[657] , \data_buffer[656] , 
            \data_buffer[652] , \data_buffer[651] , \data_buffer[650] , 
            \data_buffer[649] , \data_buffer[648] , \data_buffer[644] , 
            \data_buffer[643] , \data_buffer[642] , \data_buffer[641] , 
            \data_buffer[640] , \data_buffer[636] , \data_buffer[635] , 
            \data_buffer[634] , \data_buffer[633] , \data_buffer[632] , 
            \data_buffer[628] , \data_buffer[627] , \data_buffer[626] , 
            \data_buffer[625] , \data_buffer[624] , \data_buffer[620] , 
            \data_buffer[619] , \data_buffer[618] , \data_buffer[617] , 
            \data_buffer[616] , \data_buffer[612] , \data_buffer[611] , 
            \data_buffer[610] , \data_buffer[609] , \data_buffer[608] , 
            \data_buffer[604] , \data_buffer[603] , \data_buffer[602] , 
            \data_buffer[601] , \data_buffer[600] , \data_buffer[596] , 
            \data_buffer[595] , \data_buffer[594] , \data_buffer[593] , 
            \data_buffer[592] , \data_buffer[588] , \data_buffer[587] , 
            \data_buffer[586] , \data_buffer[585] , \data_buffer[584] , 
            \data_buffer[580] , \data_buffer[579] , \data_buffer[578] , 
            \data_buffer[577] , \data_buffer[576] , \data_buffer[572] , 
            \data_buffer[571] , \data_buffer[570] , \data_buffer[569] , 
            \data_buffer[568] , \data_buffer[564] , \data_buffer[563] , 
            \data_buffer[562] , \data_buffer[561] , \data_buffer[560] , 
            \data_buffer[556] , \data_buffer[555] , \data_buffer[554] , 
            \data_buffer[553] , \data_buffer[552] , \data_buffer[548] , 
            \data_buffer[547] , \data_buffer[546] , \data_buffer[545] , 
            \data_buffer[544] , \data_buffer[540] , \data_buffer[539] , 
            \data_buffer[538] , \data_buffer[537] , \data_buffer[536] , 
            \data_buffer[532] , \data_buffer[531] , \data_buffer[530] , 
            \data_buffer[529] , \data_buffer[528] , \data_buffer[524] , 
            \data_buffer[523] , \data_buffer[522] , \data_buffer[521] , 
            \data_buffer[520] , \data_buffer[516] , \data_buffer[515] , 
            \data_buffer[514] , \data_buffer[513] , \data_buffer[512] , 
            \data_buffer[508] , \data_buffer[507] , \data_buffer[506] , 
            \data_buffer[505] , \data_buffer[504] , \data_buffer[500] , 
            \data_buffer[499] , \data_buffer[498] , \data_buffer[497] , 
            \data_buffer[496] , \data_buffer[492] , \data_buffer[491] , 
            \data_buffer[490] , \data_buffer[489] , \data_buffer[488] , 
            \data_buffer[484] , \data_buffer[483] , \data_buffer[482] , 
            \data_buffer[481] , \data_buffer[480] , \data_buffer[476] , 
            \data_buffer[475] , \data_buffer[474] , \data_buffer[473] , 
            \data_buffer[472] , \data_buffer[468] , \data_buffer[467] , 
            \data_buffer[466] , \data_buffer[465] , \data_buffer[464] , 
            \data_buffer[460] , \data_buffer[459] , \data_buffer[458] , 
            \data_buffer[457] , \data_buffer[456] , \data_buffer[452] , 
            \data_buffer[451] , \data_buffer[450] , \data_buffer[449] , 
            \data_buffer[448] , \data_buffer[444] , \data_buffer[443] , 
            \data_buffer[442] , \data_buffer[441] , \data_buffer[440] , 
            \data_buffer[436] , \data_buffer[435] , \data_buffer[434] , 
            \data_buffer[433] , \data_buffer[426] , \data_buffer[425] , 
            \data_buffer[418] , \data_buffer[417] , \data_buffer[416] , 
            \data_buffer[412] , \data_buffer[411] , \data_buffer[410] , 
            \data_buffer[409] , \data_buffer[408] , \data_buffer[404] , 
            \data_buffer[403] , \data_buffer[402] , \data_buffer[401] , 
            \data_buffer[400] , \data_buffer[396] , \data_buffer[395] , 
            \data_buffer[394] , \data_buffer[393] , \data_buffer[392] , 
            \data_buffer[388] , \data_buffer[387] , \data_buffer[386] , 
            \data_buffer[385] , \data_buffer[384] , \data_buffer[380] , 
            \data_buffer[379] , \data_buffer[378] , \data_buffer[377] , 
            \data_buffer[376] , \data_buffer[372] , \data_buffer[371] , 
            \data_buffer[370] , \data_buffer[369] , \data_buffer[368] , 
            \data_buffer[364] , \data_buffer[363] , \data_buffer[362] , 
            \data_buffer[361] , \data_buffer[360] , \data_buffer[356] , 
            \data_buffer[355] , \data_buffer[354] , \data_buffer[353] , 
            \data_buffer[352] , \data_buffer[348] , \data_buffer[347] , 
            \data_buffer[346] , \data_buffer[345] , \data_buffer[344] , 
            \data_buffer[340] , \data_buffer[339] , \data_buffer[338] , 
            \data_buffer[337] , \data_buffer[336] , \data_buffer[332] , 
            \data_buffer[331] , \data_buffer[330] , \data_buffer[329] , 
            \data_buffer[328] , \data_buffer[324] , \data_buffer[323] , 
            \data_buffer[322] , \data_buffer[321] , \data_buffer[320] , 
            \data_buffer[316] , \data_buffer[315] , \data_buffer[314] , 
            \data_buffer[313] , \data_buffer[312] , \data_buffer[308] , 
            \data_buffer[307] , \data_buffer[306] , \data_buffer[305] , 
            \data_buffer[304] , \data_buffer[300] , \data_buffer[299] , 
            \data_buffer[298] , \data_buffer[297] , \data_buffer[296] , 
            \data_buffer[292] , \data_buffer[291] , \data_buffer[290] , 
            \data_buffer[289] , \data_buffer[288] , \data_buffer[284] , 
            \data_buffer[283] , \data_buffer[282] , \data_buffer[281] , 
            \data_buffer[280] , \data_buffer[276] , \data_buffer[275] , 
            \data_buffer[274] , \data_buffer[273] , \data_buffer[272] , 
            \data_buffer[268] , \data_buffer[267] , \data_buffer[266] , 
            \data_buffer[265] , \data_buffer[264] , \data_buffer[260] , 
            \data_buffer[259] , \data_buffer[258] , \data_buffer[257] , 
            \data_buffer[256] , \data_buffer[252] , \data_buffer[251] , 
            \data_buffer[250] , \data_buffer[249] , \data_buffer[248] , 
            \data_buffer[244] , \data_buffer[243] , \data_buffer[242] , 
            \data_buffer[241] , \data_buffer[240] , \data_buffer[236] , 
            \data_buffer[235] , \data_buffer[234] , \data_buffer[233] , 
            \data_buffer[232] , \data_buffer[228] , \data_buffer[227] , 
            \data_buffer[226] , \data_buffer[225] , \data_buffer[224] , 
            \data_buffer[220] , \data_buffer[219] , \data_buffer[218] , 
            \data_buffer[217] , n26793, \data_buffer[216] , \data_buffer[212] , 
            \data_buffer[211] , \data_buffer[210] , \data_buffer[209] , 
            \data_buffer[208] , \data_buffer[204] , \data_buffer[203] , 
            \data_buffer[202] , \data_buffer[201] , \data_buffer[200] , 
            \data_buffer[196] , \data_buffer[195] , \data_buffer[194] , 
            \data_buffer[193] , \data_buffer[192] , \data_buffer[188] , 
            \data_buffer[187] , \data_buffer[178] , \data_buffer[170] , 
            \data_buffer[179] , \data_buffer[171] , \data_buffer[180] , 
            \data_buffer[172] , \data_buffer[184] , \data_buffer[176] , 
            \data_buffer[185] , \data_buffer[177] , \data_buffer[186] , 
            \data_buffer[169] , \data_buffer[168] , \data_buffer[164] , 
            \data_buffer[163] , \data_buffer[162] , \data_buffer[161] , 
            \data_buffer[160] , \data_buffer[156] , \data_buffer[155] , 
            \data_buffer[154] , \data_buffer[153] , \data_buffer[152] , 
            \data_buffer[148] , \data_buffer[147] , \data_buffer[146] , 
            \data_buffer[145] , \data_buffer[144] , \data_buffer[140] , 
            \data_buffer[139] , \data_buffer[138] , \data_buffer[137] , 
            \data_buffer[136] , \data_buffer[132] , \data_buffer[131] , 
            \data_buffer[130] , \data_buffer[129] , \data_buffer[128] , 
            \data_buffer[124] , \data_buffer[123] , \data_buffer[122] , 
            \data_buffer[121] , \data_buffer[120] , \data_buffer[116] , 
            \data_buffer[115] , \data_buffer[114] , \data_buffer[113] , 
            \data_buffer[112] , \data_buffer[108] , \data_buffer[107] , 
            \data_buffer[106] , \data_buffer[105] , \data_buffer[104] , 
            \data_buffer[100] , \data_buffer[99] , \data_buffer[98] , 
            \data_buffer[97] , \data_buffer[96] , \data_buffer[92] , \data_buffer[91] , 
            \data_buffer[90] , \data_buffer[89] , \data_buffer[88] , \data_buffer[84] , 
            \data_buffer[83] , \data_buffer[82] , \data_buffer[81] , \data_buffer[80] , 
            \data_buffer[76] , \data_buffer[75] , \data_buffer[74] , \data_buffer[73] , 
            data_length, clk_c_enable_1399, \data_buffer[72] , \data_buffer[68] , 
            \data_buffer[67] , \data_buffer[66] , \data_buffer[65] , \data_buffer[64] , 
            \data_buffer[60] , \data_buffer[59] , \data_buffer[58] , \data_buffer[57] , 
            \data_buffer[56] , \data_buffer[52] , \data_buffer[51] , \data_buffer[50] , 
            \data_buffer[49] , \data_buffer[48] , \data_buffer[44] , \data_buffer[43] , 
            \data_buffer[42] , \data_buffer[41] , \data_buffer[40] , \data_buffer[36] , 
            \data_buffer[35] , \data_buffer[34] , \data_buffer[33] , \data_buffer[32] , 
            \data_buffer[28] , \data_buffer[27] , \data_buffer[26] , \data_buffer[25] , 
            \data_buffer[24] , \data_buffer[20] , \data_buffer[19] , \data_buffer[18] , 
            \data_buffer[17] , \data_buffer[16] , \data_buffer[12] , \data_buffer[11] , 
            \data_buffer[10] , \data_buffer[9] , \data_buffer[8] , \data_buffer[4] , 
            \data_buffer[3] , \data_buffer[2] , \data_buffer[1] , flag, 
            GND_net, \tamp_data[0] , \tamp_data[4] , \tamp_data[1] , 
            \tamp_data[5] , \tamp_data[2] , \tamp_data[6] , \tamp_data[3] , 
            \tamp_data[7] , \tamp_data[9] , \tamp_data[8] , n15, ready, 
            rs232_tx_c, rs232_rx_c) /* synthesis syn_module_defined=1 */ ;
    output \data_buffer[432] ;
    input clk_c;
    input clk_c_enable_659;
    output \data_buffer[424] ;
    output \data_buffer[0] ;
    output \data_buffer[956] ;
    output \data_buffer[948] ;
    output \data_buffer[955] ;
    output \data_buffer[947] ;
    output \data_buffer[954] ;
    output \data_buffer[946] ;
    output \data_buffer[953] ;
    output \data_buffer[945] ;
    output \data_buffer[952] ;
    output \data_buffer[944] ;
    output \data_buffer[940] ;
    output \data_buffer[939] ;
    output \data_buffer[938] ;
    output \data_buffer[937] ;
    output \data_buffer[936] ;
    output \data_buffer[932] ;
    output \data_buffer[931] ;
    output \data_buffer[930] ;
    output \data_buffer[929] ;
    output \data_buffer[928] ;
    output \data_buffer[924] ;
    output \data_buffer[923] ;
    output \data_buffer[922] ;
    output \data_buffer[921] ;
    output \data_buffer[920] ;
    output \data_buffer[916] ;
    output \data_buffer[915] ;
    output \data_buffer[914] ;
    output \data_buffer[913] ;
    output \data_buffer[912] ;
    output \data_buffer[908] ;
    output \data_buffer[907] ;
    output \data_buffer[906] ;
    output \data_buffer[905] ;
    output \data_buffer[904] ;
    output \data_buffer[900] ;
    output \data_buffer[899] ;
    output \data_buffer[898] ;
    output \data_buffer[897] ;
    output \data_buffer[896] ;
    output \data_buffer[892] ;
    output \data_buffer[891] ;
    output \data_buffer[428] ;
    output \data_buffer[420] ;
    output \data_buffer[427] ;
    output \data_buffer[419] ;
    output \data_buffer[890] ;
    output \data_buffer[889] ;
    output \data_buffer[888] ;
    output \data_buffer[884] ;
    output \data_buffer[883] ;
    output \data_buffer[882] ;
    output \data_buffer[881] ;
    output \data_buffer[880] ;
    output \data_buffer[876] ;
    output \data_buffer[875] ;
    output \data_buffer[874] ;
    output \data_buffer[873] ;
    output \data_buffer[872] ;
    output \data_buffer[868] ;
    output \data_buffer[867] ;
    output \data_buffer[866] ;
    output \data_buffer[865] ;
    output \data_buffer[864] ;
    output \data_buffer[860] ;
    output \data_buffer[859] ;
    output \data_buffer[858] ;
    output \data_buffer[857] ;
    output \data_buffer[856] ;
    output \data_buffer[852] ;
    output \data_buffer[851] ;
    output \data_buffer[850] ;
    output \data_buffer[849] ;
    output \data_buffer[848] ;
    output \data_buffer[844] ;
    output \data_buffer[843] ;
    output \data_buffer[842] ;
    output \data_buffer[841] ;
    output \data_buffer[840] ;
    output \data_buffer[836] ;
    output \data_buffer[835] ;
    output \data_buffer[834] ;
    output \data_buffer[833] ;
    output \data_buffer[832] ;
    output \data_buffer[828] ;
    output \data_buffer[827] ;
    output \data_buffer[826] ;
    output \data_buffer[825] ;
    output \data_buffer[824] ;
    output \data_buffer[820] ;
    output \data_buffer[819] ;
    output \data_buffer[818] ;
    output \data_buffer[817] ;
    output \data_buffer[816] ;
    output \data_buffer[812] ;
    output \data_buffer[811] ;
    output \data_buffer[810] ;
    output \data_buffer[809] ;
    output \data_buffer[808] ;
    output \data_buffer[804] ;
    output \data_buffer[803] ;
    output \data_buffer[802] ;
    output \data_buffer[801] ;
    output \data_buffer[800] ;
    output \data_buffer[796] ;
    output \data_buffer[795] ;
    output \data_buffer[794] ;
    output \data_buffer[793] ;
    output \data_buffer[792] ;
    input n26780;
    output \data_buffer[788] ;
    output \data_buffer[787] ;
    output \data_buffer[786] ;
    output \data_buffer[785] ;
    output \data_buffer[784] ;
    output \data_buffer[780] ;
    output \data_buffer[779] ;
    output \data_buffer[778] ;
    output \data_buffer[777] ;
    output \data_buffer[776] ;
    output \data_buffer[772] ;
    output \data_buffer[771] ;
    output \data_buffer[770] ;
    output \data_buffer[769] ;
    output \data_buffer[768] ;
    output \data_buffer[764] ;
    output \data_buffer[763] ;
    output \data_buffer[762] ;
    output \data_buffer[761] ;
    output \data_buffer[760] ;
    output \data_buffer[756] ;
    output \data_buffer[755] ;
    output \data_buffer[754] ;
    output \data_buffer[753] ;
    output \data_buffer[752] ;
    output \data_buffer[748] ;
    output \data_buffer[747] ;
    output \data_buffer[746] ;
    output \data_buffer[745] ;
    output \data_buffer[744] ;
    output \data_buffer[740] ;
    output \data_buffer[739] ;
    output \data_buffer[738] ;
    output \data_buffer[737] ;
    output \data_buffer[736] ;
    output \data_buffer[732] ;
    output \data_buffer[731] ;
    output \data_buffer[730] ;
    output \data_buffer[729] ;
    output \data_buffer[728] ;
    output \data_buffer[724] ;
    output \data_buffer[723] ;
    output \data_buffer[722] ;
    output \data_buffer[721] ;
    output \data_buffer[720] ;
    output \data_buffer[716] ;
    output \data_buffer[715] ;
    output \data_buffer[714] ;
    output \data_buffer[713] ;
    output \data_buffer[712] ;
    output \data_buffer[708] ;
    output \data_buffer[707] ;
    output \data_buffer[706] ;
    output \data_buffer[705] ;
    output \data_buffer[704] ;
    output \data_buffer[700] ;
    output \data_buffer[699] ;
    output \data_buffer[698] ;
    output \data_buffer[697] ;
    output \data_buffer[696] ;
    output \data_buffer[692] ;
    output \data_buffer[691] ;
    output \data_buffer[690] ;
    output \data_buffer[689] ;
    output \data_buffer[688] ;
    output \data_buffer[684] ;
    output \data_buffer[683] ;
    output \data_buffer[682] ;
    output \data_buffer[681] ;
    output \data_buffer[680] ;
    output \data_buffer[676] ;
    output \data_buffer[675] ;
    output \data_buffer[674] ;
    output \data_buffer[673] ;
    output \data_buffer[672] ;
    output \data_buffer[668] ;
    output \data_buffer[667] ;
    output \data_buffer[666] ;
    output \data_buffer[665] ;
    output \data_buffer[664] ;
    output \data_buffer[660] ;
    output \data_buffer[659] ;
    output \data_buffer[658] ;
    output \data_buffer[657] ;
    output \data_buffer[656] ;
    output \data_buffer[652] ;
    output \data_buffer[651] ;
    output \data_buffer[650] ;
    output \data_buffer[649] ;
    output \data_buffer[648] ;
    output \data_buffer[644] ;
    output \data_buffer[643] ;
    output \data_buffer[642] ;
    output \data_buffer[641] ;
    output \data_buffer[640] ;
    output \data_buffer[636] ;
    output \data_buffer[635] ;
    output \data_buffer[634] ;
    output \data_buffer[633] ;
    output \data_buffer[632] ;
    output \data_buffer[628] ;
    output \data_buffer[627] ;
    output \data_buffer[626] ;
    output \data_buffer[625] ;
    output \data_buffer[624] ;
    output \data_buffer[620] ;
    output \data_buffer[619] ;
    output \data_buffer[618] ;
    output \data_buffer[617] ;
    output \data_buffer[616] ;
    output \data_buffer[612] ;
    output \data_buffer[611] ;
    output \data_buffer[610] ;
    output \data_buffer[609] ;
    output \data_buffer[608] ;
    output \data_buffer[604] ;
    output \data_buffer[603] ;
    output \data_buffer[602] ;
    output \data_buffer[601] ;
    output \data_buffer[600] ;
    output \data_buffer[596] ;
    output \data_buffer[595] ;
    output \data_buffer[594] ;
    output \data_buffer[593] ;
    output \data_buffer[592] ;
    output \data_buffer[588] ;
    output \data_buffer[587] ;
    output \data_buffer[586] ;
    output \data_buffer[585] ;
    output \data_buffer[584] ;
    output \data_buffer[580] ;
    output \data_buffer[579] ;
    output \data_buffer[578] ;
    output \data_buffer[577] ;
    output \data_buffer[576] ;
    output \data_buffer[572] ;
    output \data_buffer[571] ;
    output \data_buffer[570] ;
    output \data_buffer[569] ;
    output \data_buffer[568] ;
    output \data_buffer[564] ;
    output \data_buffer[563] ;
    output \data_buffer[562] ;
    output \data_buffer[561] ;
    output \data_buffer[560] ;
    output \data_buffer[556] ;
    output \data_buffer[555] ;
    output \data_buffer[554] ;
    output \data_buffer[553] ;
    output \data_buffer[552] ;
    output \data_buffer[548] ;
    output \data_buffer[547] ;
    output \data_buffer[546] ;
    output \data_buffer[545] ;
    output \data_buffer[544] ;
    output \data_buffer[540] ;
    output \data_buffer[539] ;
    output \data_buffer[538] ;
    output \data_buffer[537] ;
    output \data_buffer[536] ;
    output \data_buffer[532] ;
    output \data_buffer[531] ;
    output \data_buffer[530] ;
    output \data_buffer[529] ;
    output \data_buffer[528] ;
    output \data_buffer[524] ;
    output \data_buffer[523] ;
    output \data_buffer[522] ;
    output \data_buffer[521] ;
    output \data_buffer[520] ;
    output \data_buffer[516] ;
    output \data_buffer[515] ;
    output \data_buffer[514] ;
    output \data_buffer[513] ;
    output \data_buffer[512] ;
    output \data_buffer[508] ;
    output \data_buffer[507] ;
    output \data_buffer[506] ;
    output \data_buffer[505] ;
    output \data_buffer[504] ;
    output \data_buffer[500] ;
    output \data_buffer[499] ;
    output \data_buffer[498] ;
    output \data_buffer[497] ;
    output \data_buffer[496] ;
    output \data_buffer[492] ;
    output \data_buffer[491] ;
    output \data_buffer[490] ;
    output \data_buffer[489] ;
    output \data_buffer[488] ;
    output \data_buffer[484] ;
    output \data_buffer[483] ;
    output \data_buffer[482] ;
    output \data_buffer[481] ;
    output \data_buffer[480] ;
    output \data_buffer[476] ;
    output \data_buffer[475] ;
    output \data_buffer[474] ;
    output \data_buffer[473] ;
    output \data_buffer[472] ;
    output \data_buffer[468] ;
    output \data_buffer[467] ;
    output \data_buffer[466] ;
    output \data_buffer[465] ;
    output \data_buffer[464] ;
    output \data_buffer[460] ;
    output \data_buffer[459] ;
    output \data_buffer[458] ;
    output \data_buffer[457] ;
    output \data_buffer[456] ;
    output \data_buffer[452] ;
    output \data_buffer[451] ;
    output \data_buffer[450] ;
    output \data_buffer[449] ;
    output \data_buffer[448] ;
    output \data_buffer[444] ;
    output \data_buffer[443] ;
    output \data_buffer[442] ;
    output \data_buffer[441] ;
    output \data_buffer[440] ;
    output \data_buffer[436] ;
    output \data_buffer[435] ;
    output \data_buffer[434] ;
    output \data_buffer[433] ;
    output \data_buffer[426] ;
    output \data_buffer[425] ;
    output \data_buffer[418] ;
    output \data_buffer[417] ;
    output \data_buffer[416] ;
    output \data_buffer[412] ;
    output \data_buffer[411] ;
    output \data_buffer[410] ;
    output \data_buffer[409] ;
    output \data_buffer[408] ;
    output \data_buffer[404] ;
    output \data_buffer[403] ;
    output \data_buffer[402] ;
    output \data_buffer[401] ;
    output \data_buffer[400] ;
    output \data_buffer[396] ;
    output \data_buffer[395] ;
    output \data_buffer[394] ;
    output \data_buffer[393] ;
    output \data_buffer[392] ;
    output \data_buffer[388] ;
    output \data_buffer[387] ;
    output \data_buffer[386] ;
    output \data_buffer[385] ;
    output \data_buffer[384] ;
    output \data_buffer[380] ;
    output \data_buffer[379] ;
    output \data_buffer[378] ;
    output \data_buffer[377] ;
    output \data_buffer[376] ;
    output \data_buffer[372] ;
    output \data_buffer[371] ;
    output \data_buffer[370] ;
    output \data_buffer[369] ;
    output \data_buffer[368] ;
    output \data_buffer[364] ;
    output \data_buffer[363] ;
    output \data_buffer[362] ;
    output \data_buffer[361] ;
    output \data_buffer[360] ;
    output \data_buffer[356] ;
    output \data_buffer[355] ;
    output \data_buffer[354] ;
    output \data_buffer[353] ;
    output \data_buffer[352] ;
    output \data_buffer[348] ;
    output \data_buffer[347] ;
    output \data_buffer[346] ;
    output \data_buffer[345] ;
    output \data_buffer[344] ;
    output \data_buffer[340] ;
    output \data_buffer[339] ;
    output \data_buffer[338] ;
    output \data_buffer[337] ;
    output \data_buffer[336] ;
    output \data_buffer[332] ;
    output \data_buffer[331] ;
    output \data_buffer[330] ;
    output \data_buffer[329] ;
    output \data_buffer[328] ;
    output \data_buffer[324] ;
    output \data_buffer[323] ;
    output \data_buffer[322] ;
    output \data_buffer[321] ;
    output \data_buffer[320] ;
    output \data_buffer[316] ;
    output \data_buffer[315] ;
    output \data_buffer[314] ;
    output \data_buffer[313] ;
    output \data_buffer[312] ;
    output \data_buffer[308] ;
    output \data_buffer[307] ;
    output \data_buffer[306] ;
    output \data_buffer[305] ;
    output \data_buffer[304] ;
    output \data_buffer[300] ;
    output \data_buffer[299] ;
    output \data_buffer[298] ;
    output \data_buffer[297] ;
    output \data_buffer[296] ;
    output \data_buffer[292] ;
    output \data_buffer[291] ;
    output \data_buffer[290] ;
    output \data_buffer[289] ;
    output \data_buffer[288] ;
    output \data_buffer[284] ;
    output \data_buffer[283] ;
    output \data_buffer[282] ;
    output \data_buffer[281] ;
    output \data_buffer[280] ;
    output \data_buffer[276] ;
    output \data_buffer[275] ;
    output \data_buffer[274] ;
    output \data_buffer[273] ;
    output \data_buffer[272] ;
    output \data_buffer[268] ;
    output \data_buffer[267] ;
    output \data_buffer[266] ;
    output \data_buffer[265] ;
    output \data_buffer[264] ;
    output \data_buffer[260] ;
    output \data_buffer[259] ;
    output \data_buffer[258] ;
    output \data_buffer[257] ;
    output \data_buffer[256] ;
    output \data_buffer[252] ;
    output \data_buffer[251] ;
    output \data_buffer[250] ;
    output \data_buffer[249] ;
    output \data_buffer[248] ;
    output \data_buffer[244] ;
    output \data_buffer[243] ;
    output \data_buffer[242] ;
    output \data_buffer[241] ;
    output \data_buffer[240] ;
    output \data_buffer[236] ;
    output \data_buffer[235] ;
    output \data_buffer[234] ;
    output \data_buffer[233] ;
    output \data_buffer[232] ;
    output \data_buffer[228] ;
    output \data_buffer[227] ;
    output \data_buffer[226] ;
    output \data_buffer[225] ;
    output \data_buffer[224] ;
    output \data_buffer[220] ;
    output \data_buffer[219] ;
    output \data_buffer[218] ;
    output \data_buffer[217] ;
    output n26793;
    output \data_buffer[216] ;
    output \data_buffer[212] ;
    output \data_buffer[211] ;
    output \data_buffer[210] ;
    output \data_buffer[209] ;
    output \data_buffer[208] ;
    output \data_buffer[204] ;
    output \data_buffer[203] ;
    output \data_buffer[202] ;
    output \data_buffer[201] ;
    output \data_buffer[200] ;
    output \data_buffer[196] ;
    output \data_buffer[195] ;
    output \data_buffer[194] ;
    output \data_buffer[193] ;
    output \data_buffer[192] ;
    output \data_buffer[188] ;
    output \data_buffer[187] ;
    output \data_buffer[178] ;
    output \data_buffer[170] ;
    output \data_buffer[179] ;
    output \data_buffer[171] ;
    output \data_buffer[180] ;
    output \data_buffer[172] ;
    output \data_buffer[184] ;
    output \data_buffer[176] ;
    output \data_buffer[185] ;
    output \data_buffer[177] ;
    output \data_buffer[186] ;
    output \data_buffer[169] ;
    output \data_buffer[168] ;
    output \data_buffer[164] ;
    output \data_buffer[163] ;
    output \data_buffer[162] ;
    output \data_buffer[161] ;
    output \data_buffer[160] ;
    output \data_buffer[156] ;
    output \data_buffer[155] ;
    output \data_buffer[154] ;
    output \data_buffer[153] ;
    output \data_buffer[152] ;
    output \data_buffer[148] ;
    output \data_buffer[147] ;
    output \data_buffer[146] ;
    output \data_buffer[145] ;
    output \data_buffer[144] ;
    output \data_buffer[140] ;
    output \data_buffer[139] ;
    output \data_buffer[138] ;
    output \data_buffer[137] ;
    output \data_buffer[136] ;
    output \data_buffer[132] ;
    output \data_buffer[131] ;
    output \data_buffer[130] ;
    output \data_buffer[129] ;
    output \data_buffer[128] ;
    output \data_buffer[124] ;
    output \data_buffer[123] ;
    output \data_buffer[122] ;
    output \data_buffer[121] ;
    output \data_buffer[120] ;
    output \data_buffer[116] ;
    output \data_buffer[115] ;
    output \data_buffer[114] ;
    output \data_buffer[113] ;
    output \data_buffer[112] ;
    output \data_buffer[108] ;
    output \data_buffer[107] ;
    output \data_buffer[106] ;
    output \data_buffer[105] ;
    output \data_buffer[104] ;
    output \data_buffer[100] ;
    output \data_buffer[99] ;
    output \data_buffer[98] ;
    output \data_buffer[97] ;
    output \data_buffer[96] ;
    output \data_buffer[92] ;
    output \data_buffer[91] ;
    output \data_buffer[90] ;
    output \data_buffer[89] ;
    output \data_buffer[88] ;
    output \data_buffer[84] ;
    output \data_buffer[83] ;
    output \data_buffer[82] ;
    output \data_buffer[81] ;
    output \data_buffer[80] ;
    output \data_buffer[76] ;
    output \data_buffer[75] ;
    output \data_buffer[74] ;
    output \data_buffer[73] ;
    output [9:0]data_length;
    input clk_c_enable_1399;
    output \data_buffer[72] ;
    output \data_buffer[68] ;
    output \data_buffer[67] ;
    output \data_buffer[66] ;
    output \data_buffer[65] ;
    output \data_buffer[64] ;
    output \data_buffer[60] ;
    output \data_buffer[59] ;
    output \data_buffer[58] ;
    output \data_buffer[57] ;
    output \data_buffer[56] ;
    output \data_buffer[52] ;
    output \data_buffer[51] ;
    output \data_buffer[50] ;
    output \data_buffer[49] ;
    output \data_buffer[48] ;
    output \data_buffer[44] ;
    output \data_buffer[43] ;
    output \data_buffer[42] ;
    output \data_buffer[41] ;
    output \data_buffer[40] ;
    output \data_buffer[36] ;
    output \data_buffer[35] ;
    output \data_buffer[34] ;
    output \data_buffer[33] ;
    output \data_buffer[32] ;
    output \data_buffer[28] ;
    output \data_buffer[27] ;
    output \data_buffer[26] ;
    output \data_buffer[25] ;
    output \data_buffer[24] ;
    output \data_buffer[20] ;
    output \data_buffer[19] ;
    output \data_buffer[18] ;
    output \data_buffer[17] ;
    output \data_buffer[16] ;
    output \data_buffer[12] ;
    output \data_buffer[11] ;
    output \data_buffer[10] ;
    output \data_buffer[9] ;
    output \data_buffer[8] ;
    output \data_buffer[4] ;
    output \data_buffer[3] ;
    output \data_buffer[2] ;
    output \data_buffer[1] ;
    input flag;
    input GND_net;
    input \tamp_data[0] ;
    input \tamp_data[4] ;
    input \tamp_data[1] ;
    input \tamp_data[5] ;
    input \tamp_data[2] ;
    input \tamp_data[6] ;
    input \tamp_data[3] ;
    input \tamp_data[7] ;
    input \tamp_data[9] ;
    input \tamp_data[8] ;
    output n15;
    output ready;
    output rs232_tx_c;
    input rs232_rx_c;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // g:/fpga/mxo2/system/project/system_top.v(2[15:18])
    
    wire n26798, n26802;
    wire [7:0]rx_data;   // g:/fpga/mxo2/system/project/uart_top.v(20[14:21])
    
    wire n26804, rx_done;
    wire [1:0]tx_data_length;   // g:/fpga/mxo2/system/project/uart_top.v(21[25:39])
    wire [1:0]tx_data_length_1__N_1866;
    
    wire bps_en_tx1, bps_en_tx0, bps_en_tx2;
    wire [7:0]tx_data;   // g:/fpga/mxo2/system/project/uart_top.v(52[25:32])
    
    wire clk_c_enable_1418;
    wire [7:0]tx_data_7__N_1868;
    
    wire bps_en_N_2978, tx_en, bps_en_tx, n26803, n26797, rx_done_N_2858, 
        n26794, n26799, n26805, n26801, n26800, n26795, n26796;
    wire [9:0]n78;
    
    wire tx_done, n9394, n12084, n20509, n20508, n20507, n20506, 
        n20505, n9, n23801, bps_clk_tx, bps_en_rx, bps_clk_rx;
    
    FD1P3IX data_buffer__i432 (.D(\data_buffer[424] ), .SP(clk_c_enable_659), 
            .CD(n26798), .CK(clk_c), .Q(\data_buffer[432] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i432.GSR = "ENABLED";
    FD1P3IX data_buffer__i0 (.D(rx_data[0]), .SP(clk_c_enable_659), .CD(n26802), 
            .CK(clk_c), .Q(\data_buffer[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i0.GSR = "ENABLED";
    FD1P3IX data_buffer__i956 (.D(\data_buffer[948] ), .SP(clk_c_enable_659), 
            .CD(n26804), .CK(clk_c), .Q(\data_buffer[956] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i956.GSR = "ENABLED";
    FD1P3IX data_buffer__i955 (.D(\data_buffer[947] ), .SP(clk_c_enable_659), 
            .CD(rx_done), .CK(clk_c), .Q(\data_buffer[955] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i955.GSR = "ENABLED";
    FD1P3IX data_buffer__i954 (.D(\data_buffer[946] ), .SP(clk_c_enable_659), 
            .CD(n26804), .CK(clk_c), .Q(\data_buffer[954] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i954.GSR = "ENABLED";
    FD1P3IX data_buffer__i953 (.D(\data_buffer[945] ), .SP(clk_c_enable_659), 
            .CD(rx_done), .CK(clk_c), .Q(\data_buffer[953] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i953.GSR = "ENABLED";
    FD1P3IX data_buffer__i952 (.D(\data_buffer[944] ), .SP(clk_c_enable_659), 
            .CD(rx_done), .CK(clk_c), .Q(\data_buffer[952] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i952.GSR = "ENABLED";
    FD1P3IX data_buffer__i948 (.D(\data_buffer[940] ), .SP(clk_c_enable_659), 
            .CD(n26804), .CK(clk_c), .Q(\data_buffer[948] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i948.GSR = "ENABLED";
    FD1P3IX data_buffer__i947 (.D(\data_buffer[939] ), .SP(clk_c_enable_659), 
            .CD(rx_done), .CK(clk_c), .Q(\data_buffer[947] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i947.GSR = "ENABLED";
    FD1P3IX data_buffer__i946 (.D(\data_buffer[938] ), .SP(clk_c_enable_659), 
            .CD(n26802), .CK(clk_c), .Q(\data_buffer[946] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i946.GSR = "ENABLED";
    FD1P3IX data_buffer__i945 (.D(\data_buffer[937] ), .SP(clk_c_enable_659), 
            .CD(rx_done), .CK(clk_c), .Q(\data_buffer[945] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i945.GSR = "ENABLED";
    FD1P3IX data_buffer__i944 (.D(\data_buffer[936] ), .SP(clk_c_enable_659), 
            .CD(n26798), .CK(clk_c), .Q(\data_buffer[944] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i944.GSR = "ENABLED";
    FD1S3AX tx_data_length_i0 (.D(tx_data_length_1__N_1866[0]), .CK(clk_c), 
            .Q(tx_data_length[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(46[10] 49[49])
    defparam tx_data_length_i0.GSR = "ENABLED";
    FD1S3AX bps_en_tx1_57 (.D(bps_en_tx0), .CK(clk_c), .Q(bps_en_tx1)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(32[11] 36[5])
    defparam bps_en_tx1_57.GSR = "ENABLED";
    FD1S3AX bps_en_tx2_58 (.D(bps_en_tx1), .CK(clk_c), .Q(bps_en_tx2)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(32[11] 36[5])
    defparam bps_en_tx2_58.GSR = "ENABLED";
    FD1P3AX tx_data_i0 (.D(tx_data_7__N_1868[0]), .SP(clk_c_enable_1418), 
            .CK(clk_c), .Q(tx_data[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(56[10] 59[42])
    defparam tx_data_i0.GSR = "ENABLED";
    FD1S3AX tx_en_r_61 (.D(tx_en), .CK(clk_c), .Q(bps_en_N_2978)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(71[9:26])
    defparam tx_en_r_61.GSR = "ENABLED";
    FD1S3AX bps_en_tx0_56 (.D(bps_en_tx), .CK(clk_c), .Q(bps_en_tx0)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(32[11] 36[5])
    defparam bps_en_tx0_56.GSR = "ENABLED";
    FD1P3IX data_buffer__i940 (.D(\data_buffer[932] ), .SP(clk_c_enable_659), 
            .CD(n26802), .CK(clk_c), .Q(\data_buffer[940] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i940.GSR = "ENABLED";
    FD1P3IX data_buffer__i939 (.D(\data_buffer[931] ), .SP(clk_c_enable_659), 
            .CD(n26802), .CK(clk_c), .Q(\data_buffer[939] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i939.GSR = "ENABLED";
    FD1P3IX data_buffer__i938 (.D(\data_buffer[930] ), .SP(clk_c_enable_659), 
            .CD(rx_done), .CK(clk_c), .Q(\data_buffer[938] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i938.GSR = "ENABLED";
    FD1P3IX data_buffer__i937 (.D(\data_buffer[929] ), .SP(clk_c_enable_659), 
            .CD(n26804), .CK(clk_c), .Q(\data_buffer[937] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i937.GSR = "ENABLED";
    FD1P3IX data_buffer__i936 (.D(\data_buffer[928] ), .SP(clk_c_enable_659), 
            .CD(n26798), .CK(clk_c), .Q(\data_buffer[936] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i936.GSR = "ENABLED";
    FD1P3IX data_buffer__i932 (.D(\data_buffer[924] ), .SP(clk_c_enable_659), 
            .CD(n26798), .CK(clk_c), .Q(\data_buffer[932] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i932.GSR = "ENABLED";
    FD1P3IX data_buffer__i931 (.D(\data_buffer[923] ), .SP(clk_c_enable_659), 
            .CD(n26798), .CK(clk_c), .Q(\data_buffer[931] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i931.GSR = "ENABLED";
    FD1P3IX data_buffer__i930 (.D(\data_buffer[922] ), .SP(clk_c_enable_659), 
            .CD(rx_done), .CK(clk_c), .Q(\data_buffer[930] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i930.GSR = "ENABLED";
    FD1P3IX data_buffer__i929 (.D(\data_buffer[921] ), .SP(clk_c_enable_659), 
            .CD(n26798), .CK(clk_c), .Q(\data_buffer[929] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i929.GSR = "ENABLED";
    FD1P3IX data_buffer__i928 (.D(\data_buffer[920] ), .SP(clk_c_enable_659), 
            .CD(n26798), .CK(clk_c), .Q(\data_buffer[928] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i928.GSR = "ENABLED";
    FD1P3IX data_buffer__i924 (.D(\data_buffer[916] ), .SP(clk_c_enable_659), 
            .CD(n26802), .CK(clk_c), .Q(\data_buffer[924] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i924.GSR = "ENABLED";
    FD1P3IX data_buffer__i923 (.D(\data_buffer[915] ), .SP(clk_c_enable_659), 
            .CD(rx_done), .CK(clk_c), .Q(\data_buffer[923] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i923.GSR = "ENABLED";
    FD1P3IX data_buffer__i922 (.D(\data_buffer[914] ), .SP(clk_c_enable_659), 
            .CD(n26804), .CK(clk_c), .Q(\data_buffer[922] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i922.GSR = "ENABLED";
    FD1P3IX data_buffer__i921 (.D(\data_buffer[913] ), .SP(clk_c_enable_659), 
            .CD(n26802), .CK(clk_c), .Q(\data_buffer[921] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i921.GSR = "ENABLED";
    FD1P3IX data_buffer__i920 (.D(\data_buffer[912] ), .SP(clk_c_enable_659), 
            .CD(rx_done), .CK(clk_c), .Q(\data_buffer[920] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i920.GSR = "ENABLED";
    FD1P3IX data_buffer__i916 (.D(\data_buffer[908] ), .SP(clk_c_enable_659), 
            .CD(n26804), .CK(clk_c), .Q(\data_buffer[916] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i916.GSR = "ENABLED";
    FD1P3IX data_buffer__i915 (.D(\data_buffer[907] ), .SP(clk_c_enable_659), 
            .CD(n26802), .CK(clk_c), .Q(\data_buffer[915] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i915.GSR = "ENABLED";
    FD1P3IX data_buffer__i914 (.D(\data_buffer[906] ), .SP(clk_c_enable_659), 
            .CD(n26804), .CK(clk_c), .Q(\data_buffer[914] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i914.GSR = "ENABLED";
    FD1P3IX data_buffer__i913 (.D(\data_buffer[905] ), .SP(clk_c_enable_659), 
            .CD(n26803), .CK(clk_c), .Q(\data_buffer[913] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i913.GSR = "ENABLED";
    FD1P3IX data_buffer__i912 (.D(\data_buffer[904] ), .SP(clk_c_enable_659), 
            .CD(n26804), .CK(clk_c), .Q(\data_buffer[912] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i912.GSR = "ENABLED";
    FD1P3IX data_buffer__i908 (.D(\data_buffer[900] ), .SP(clk_c_enable_659), 
            .CD(n26803), .CK(clk_c), .Q(\data_buffer[908] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i908.GSR = "ENABLED";
    FD1P3IX data_buffer__i907 (.D(\data_buffer[899] ), .SP(clk_c_enable_659), 
            .CD(n26804), .CK(clk_c), .Q(\data_buffer[907] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i907.GSR = "ENABLED";
    FD1P3IX data_buffer__i906 (.D(\data_buffer[898] ), .SP(clk_c_enable_659), 
            .CD(n26803), .CK(clk_c), .Q(\data_buffer[906] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i906.GSR = "ENABLED";
    FD1P3IX data_buffer__i905 (.D(\data_buffer[897] ), .SP(clk_c_enable_659), 
            .CD(n26804), .CK(clk_c), .Q(\data_buffer[905] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i905.GSR = "ENABLED";
    FD1P3IX data_buffer__i904 (.D(\data_buffer[896] ), .SP(clk_c_enable_659), 
            .CD(n26804), .CK(clk_c), .Q(\data_buffer[904] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i904.GSR = "ENABLED";
    FD1P3IX data_buffer__i900 (.D(\data_buffer[892] ), .SP(clk_c_enable_659), 
            .CD(n26804), .CK(clk_c), .Q(\data_buffer[900] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i900.GSR = "ENABLED";
    FD1P3IX data_buffer__i899 (.D(\data_buffer[891] ), .SP(clk_c_enable_659), 
            .CD(n26804), .CK(clk_c), .Q(\data_buffer[899] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i899.GSR = "ENABLED";
    FD1P3IX data_buffer__i428 (.D(\data_buffer[420] ), .SP(clk_c_enable_659), 
            .CD(n26804), .CK(clk_c), .Q(\data_buffer[428] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i428.GSR = "ENABLED";
    FD1P3IX data_buffer__i427 (.D(\data_buffer[419] ), .SP(clk_c_enable_659), 
            .CD(n26804), .CK(clk_c), .Q(\data_buffer[427] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i427.GSR = "ENABLED";
    FD1P3IX data_buffer__i898 (.D(\data_buffer[890] ), .SP(clk_c_enable_659), 
            .CD(n26804), .CK(clk_c), .Q(\data_buffer[898] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i898.GSR = "ENABLED";
    FD1P3IX data_buffer__i897 (.D(\data_buffer[889] ), .SP(clk_c_enable_659), 
            .CD(n26804), .CK(clk_c), .Q(\data_buffer[897] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i897.GSR = "ENABLED";
    FD1P3IX data_buffer__i896 (.D(\data_buffer[888] ), .SP(clk_c_enable_659), 
            .CD(n26804), .CK(clk_c), .Q(\data_buffer[896] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i896.GSR = "ENABLED";
    FD1P3IX data_buffer__i892 (.D(\data_buffer[884] ), .SP(clk_c_enable_659), 
            .CD(n26804), .CK(clk_c), .Q(\data_buffer[892] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i892.GSR = "ENABLED";
    FD1P3IX data_buffer__i891 (.D(\data_buffer[883] ), .SP(clk_c_enable_659), 
            .CD(n26804), .CK(clk_c), .Q(\data_buffer[891] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i891.GSR = "ENABLED";
    FD1P3IX data_buffer__i890 (.D(\data_buffer[882] ), .SP(clk_c_enable_659), 
            .CD(n26804), .CK(clk_c), .Q(\data_buffer[890] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i890.GSR = "ENABLED";
    FD1P3IX data_buffer__i889 (.D(\data_buffer[881] ), .SP(clk_c_enable_659), 
            .CD(n26804), .CK(clk_c), .Q(\data_buffer[889] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i889.GSR = "ENABLED";
    FD1P3IX data_buffer__i888 (.D(\data_buffer[880] ), .SP(clk_c_enable_659), 
            .CD(n26804), .CK(clk_c), .Q(\data_buffer[888] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i888.GSR = "ENABLED";
    FD1P3IX data_buffer__i884 (.D(\data_buffer[876] ), .SP(clk_c_enable_659), 
            .CD(n26804), .CK(clk_c), .Q(\data_buffer[884] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i884.GSR = "ENABLED";
    FD1P3IX data_buffer__i883 (.D(\data_buffer[875] ), .SP(clk_c_enable_659), 
            .CD(n26803), .CK(clk_c), .Q(\data_buffer[883] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i883.GSR = "ENABLED";
    FD1P3IX data_buffer__i882 (.D(\data_buffer[874] ), .SP(clk_c_enable_659), 
            .CD(n26804), .CK(clk_c), .Q(\data_buffer[882] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i882.GSR = "ENABLED";
    FD1P3IX data_buffer__i881 (.D(\data_buffer[873] ), .SP(clk_c_enable_659), 
            .CD(n26803), .CK(clk_c), .Q(\data_buffer[881] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i881.GSR = "ENABLED";
    FD1P3IX data_buffer__i880 (.D(\data_buffer[872] ), .SP(clk_c_enable_659), 
            .CD(n26804), .CK(clk_c), .Q(\data_buffer[880] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i880.GSR = "ENABLED";
    FD1P3IX data_buffer__i876 (.D(\data_buffer[868] ), .SP(clk_c_enable_659), 
            .CD(n26803), .CK(clk_c), .Q(\data_buffer[876] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i876.GSR = "ENABLED";
    FD1P3IX data_buffer__i875 (.D(\data_buffer[867] ), .SP(clk_c_enable_659), 
            .CD(n26804), .CK(clk_c), .Q(\data_buffer[875] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i875.GSR = "ENABLED";
    FD1P3IX data_buffer__i874 (.D(\data_buffer[866] ), .SP(clk_c_enable_659), 
            .CD(n26803), .CK(clk_c), .Q(\data_buffer[874] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i874.GSR = "ENABLED";
    FD1P3IX data_buffer__i873 (.D(\data_buffer[865] ), .SP(clk_c_enable_659), 
            .CD(n26804), .CK(clk_c), .Q(\data_buffer[873] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i873.GSR = "ENABLED";
    FD1P3IX data_buffer__i872 (.D(\data_buffer[864] ), .SP(clk_c_enable_659), 
            .CD(n26803), .CK(clk_c), .Q(\data_buffer[872] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i872.GSR = "ENABLED";
    FD1P3IX data_buffer__i868 (.D(\data_buffer[860] ), .SP(clk_c_enable_659), 
            .CD(n26804), .CK(clk_c), .Q(\data_buffer[868] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i868.GSR = "ENABLED";
    FD1P3IX data_buffer__i867 (.D(\data_buffer[859] ), .SP(clk_c_enable_659), 
            .CD(n26803), .CK(clk_c), .Q(\data_buffer[867] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i867.GSR = "ENABLED";
    FD1P3IX data_buffer__i866 (.D(\data_buffer[858] ), .SP(clk_c_enable_659), 
            .CD(n26804), .CK(clk_c), .Q(\data_buffer[866] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i866.GSR = "ENABLED";
    FD1P3IX data_buffer__i865 (.D(\data_buffer[857] ), .SP(clk_c_enable_659), 
            .CD(n26803), .CK(clk_c), .Q(\data_buffer[865] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i865.GSR = "ENABLED";
    FD1P3IX data_buffer__i864 (.D(\data_buffer[856] ), .SP(clk_c_enable_659), 
            .CD(n26804), .CK(clk_c), .Q(\data_buffer[864] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i864.GSR = "ENABLED";
    FD1P3IX data_buffer__i860 (.D(\data_buffer[852] ), .SP(clk_c_enable_659), 
            .CD(n26798), .CK(clk_c), .Q(\data_buffer[860] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i860.GSR = "ENABLED";
    FD1P3IX data_buffer__i859 (.D(\data_buffer[851] ), .SP(clk_c_enable_659), 
            .CD(n26802), .CK(clk_c), .Q(\data_buffer[859] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i859.GSR = "ENABLED";
    FD1P3IX data_buffer__i858 (.D(\data_buffer[850] ), .SP(clk_c_enable_659), 
            .CD(n26803), .CK(clk_c), .Q(\data_buffer[858] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i858.GSR = "ENABLED";
    FD1P3IX data_buffer__i857 (.D(\data_buffer[849] ), .SP(clk_c_enable_659), 
            .CD(n26804), .CK(clk_c), .Q(\data_buffer[857] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i857.GSR = "ENABLED";
    FD1P3IX data_buffer__i856 (.D(\data_buffer[848] ), .SP(clk_c_enable_659), 
            .CD(n26802), .CK(clk_c), .Q(\data_buffer[856] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i856.GSR = "ENABLED";
    FD1P3IX data_buffer__i852 (.D(\data_buffer[844] ), .SP(clk_c_enable_659), 
            .CD(n26803), .CK(clk_c), .Q(\data_buffer[852] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i852.GSR = "ENABLED";
    FD1P3IX data_buffer__i851 (.D(\data_buffer[843] ), .SP(clk_c_enable_659), 
            .CD(n26804), .CK(clk_c), .Q(\data_buffer[851] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i851.GSR = "ENABLED";
    FD1P3IX data_buffer__i850 (.D(\data_buffer[842] ), .SP(clk_c_enable_659), 
            .CD(n26803), .CK(clk_c), .Q(\data_buffer[850] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i850.GSR = "ENABLED";
    FD1P3IX data_buffer__i849 (.D(\data_buffer[841] ), .SP(clk_c_enable_659), 
            .CD(n26802), .CK(clk_c), .Q(\data_buffer[849] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i849.GSR = "ENABLED";
    FD1P3IX data_buffer__i848 (.D(\data_buffer[840] ), .SP(clk_c_enable_659), 
            .CD(n26803), .CK(clk_c), .Q(\data_buffer[848] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i848.GSR = "ENABLED";
    FD1P3IX data_buffer__i844 (.D(\data_buffer[836] ), .SP(clk_c_enable_659), 
            .CD(n26803), .CK(clk_c), .Q(\data_buffer[844] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i844.GSR = "ENABLED";
    FD1P3IX data_buffer__i843 (.D(\data_buffer[835] ), .SP(clk_c_enable_659), 
            .CD(n26804), .CK(clk_c), .Q(\data_buffer[843] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i843.GSR = "ENABLED";
    FD1P3IX data_buffer__i842 (.D(\data_buffer[834] ), .SP(clk_c_enable_659), 
            .CD(n26802), .CK(clk_c), .Q(\data_buffer[842] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i842.GSR = "ENABLED";
    FD1P3IX data_buffer__i841 (.D(\data_buffer[833] ), .SP(clk_c_enable_659), 
            .CD(n26804), .CK(clk_c), .Q(\data_buffer[841] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i841.GSR = "ENABLED";
    FD1P3IX data_buffer__i840 (.D(\data_buffer[832] ), .SP(clk_c_enable_659), 
            .CD(n26802), .CK(clk_c), .Q(\data_buffer[840] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i840.GSR = "ENABLED";
    FD1P3IX data_buffer__i836 (.D(\data_buffer[828] ), .SP(clk_c_enable_659), 
            .CD(n26802), .CK(clk_c), .Q(\data_buffer[836] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i836.GSR = "ENABLED";
    FD1P3IX data_buffer__i835 (.D(\data_buffer[827] ), .SP(clk_c_enable_659), 
            .CD(n26804), .CK(clk_c), .Q(\data_buffer[835] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i835.GSR = "ENABLED";
    FD1P3IX data_buffer__i834 (.D(\data_buffer[826] ), .SP(clk_c_enable_659), 
            .CD(n26803), .CK(clk_c), .Q(\data_buffer[834] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i834.GSR = "ENABLED";
    FD1P3IX data_buffer__i833 (.D(\data_buffer[825] ), .SP(clk_c_enable_659), 
            .CD(n26804), .CK(clk_c), .Q(\data_buffer[833] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i833.GSR = "ENABLED";
    FD1P3IX data_buffer__i832 (.D(\data_buffer[824] ), .SP(clk_c_enable_659), 
            .CD(n26802), .CK(clk_c), .Q(\data_buffer[832] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i832.GSR = "ENABLED";
    FD1P3IX data_buffer__i828 (.D(\data_buffer[820] ), .SP(clk_c_enable_659), 
            .CD(n26802), .CK(clk_c), .Q(\data_buffer[828] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i828.GSR = "ENABLED";
    FD1P3IX data_buffer__i827 (.D(\data_buffer[819] ), .SP(clk_c_enable_659), 
            .CD(n26804), .CK(clk_c), .Q(\data_buffer[827] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i827.GSR = "ENABLED";
    FD1P3IX data_buffer__i826 (.D(\data_buffer[818] ), .SP(clk_c_enable_659), 
            .CD(n26802), .CK(clk_c), .Q(\data_buffer[826] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i826.GSR = "ENABLED";
    FD1P3IX data_buffer__i825 (.D(\data_buffer[817] ), .SP(clk_c_enable_659), 
            .CD(n26798), .CK(clk_c), .Q(\data_buffer[825] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i825.GSR = "ENABLED";
    FD1P3IX data_buffer__i824 (.D(\data_buffer[816] ), .SP(clk_c_enable_659), 
            .CD(n26798), .CK(clk_c), .Q(\data_buffer[824] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i824.GSR = "ENABLED";
    FD1P3IX data_buffer__i820 (.D(\data_buffer[812] ), .SP(clk_c_enable_659), 
            .CD(n26798), .CK(clk_c), .Q(\data_buffer[820] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i820.GSR = "ENABLED";
    FD1P3IX data_buffer__i819 (.D(\data_buffer[811] ), .SP(clk_c_enable_659), 
            .CD(n26798), .CK(clk_c), .Q(\data_buffer[819] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i819.GSR = "ENABLED";
    FD1P3IX data_buffer__i818 (.D(\data_buffer[810] ), .SP(clk_c_enable_659), 
            .CD(n26798), .CK(clk_c), .Q(\data_buffer[818] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i818.GSR = "ENABLED";
    FD1P3IX data_buffer__i817 (.D(\data_buffer[809] ), .SP(clk_c_enable_659), 
            .CD(n26803), .CK(clk_c), .Q(\data_buffer[817] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i817.GSR = "ENABLED";
    FD1P3IX data_buffer__i816 (.D(\data_buffer[808] ), .SP(clk_c_enable_659), 
            .CD(n26803), .CK(clk_c), .Q(\data_buffer[816] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i816.GSR = "ENABLED";
    FD1P3IX data_buffer__i812 (.D(\data_buffer[804] ), .SP(clk_c_enable_659), 
            .CD(n26804), .CK(clk_c), .Q(\data_buffer[812] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i812.GSR = "ENABLED";
    FD1P3IX data_buffer__i811 (.D(\data_buffer[803] ), .SP(clk_c_enable_659), 
            .CD(n26798), .CK(clk_c), .Q(\data_buffer[811] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i811.GSR = "ENABLED";
    FD1P3IX data_buffer__i810 (.D(\data_buffer[802] ), .SP(clk_c_enable_659), 
            .CD(n26798), .CK(clk_c), .Q(\data_buffer[810] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i810.GSR = "ENABLED";
    FD1P3IX data_buffer__i809 (.D(\data_buffer[801] ), .SP(clk_c_enable_659), 
            .CD(n26798), .CK(clk_c), .Q(\data_buffer[809] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i809.GSR = "ENABLED";
    FD1P3IX data_buffer__i808 (.D(\data_buffer[800] ), .SP(clk_c_enable_659), 
            .CD(n26798), .CK(clk_c), .Q(\data_buffer[808] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i808.GSR = "ENABLED";
    FD1P3IX data_buffer__i804 (.D(\data_buffer[796] ), .SP(clk_c_enable_659), 
            .CD(n26798), .CK(clk_c), .Q(\data_buffer[804] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i804.GSR = "ENABLED";
    FD1P3IX data_buffer__i803 (.D(\data_buffer[795] ), .SP(clk_c_enable_659), 
            .CD(n26802), .CK(clk_c), .Q(\data_buffer[803] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i803.GSR = "ENABLED";
    FD1P3IX data_buffer__i802 (.D(\data_buffer[794] ), .SP(clk_c_enable_659), 
            .CD(n26802), .CK(clk_c), .Q(\data_buffer[802] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i802.GSR = "ENABLED";
    FD1P3IX data_buffer__i801 (.D(\data_buffer[793] ), .SP(clk_c_enable_659), 
            .CD(n26802), .CK(clk_c), .Q(\data_buffer[801] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i801.GSR = "ENABLED";
    FD1P3IX data_buffer__i800 (.D(\data_buffer[792] ), .SP(clk_c_enable_659), 
            .CD(n26797), .CK(clk_c), .Q(\data_buffer[800] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i800.GSR = "ENABLED";
    FD1P3IX rx_done_64_rep_497 (.D(n26780), .SP(rx_done_N_2858), .CD(rx_done), 
            .CK(clk_c), .Q(n26794)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(101[10] 104[25])
    defparam rx_done_64_rep_497.GSR = "ENABLED";
    FD1P3IX data_buffer__i796 (.D(\data_buffer[788] ), .SP(clk_c_enable_659), 
            .CD(n26804), .CK(clk_c), .Q(\data_buffer[796] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i796.GSR = "ENABLED";
    FD1P3IX data_buffer__i795 (.D(\data_buffer[787] ), .SP(clk_c_enable_659), 
            .CD(n26804), .CK(clk_c), .Q(\data_buffer[795] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i795.GSR = "ENABLED";
    FD1P3IX data_buffer__i794 (.D(\data_buffer[786] ), .SP(clk_c_enable_659), 
            .CD(n26798), .CK(clk_c), .Q(\data_buffer[794] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i794.GSR = "ENABLED";
    FD1P3IX data_buffer__i793 (.D(\data_buffer[785] ), .SP(clk_c_enable_659), 
            .CD(n26799), .CK(clk_c), .Q(\data_buffer[793] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i793.GSR = "ENABLED";
    FD1P3IX data_buffer__i792 (.D(\data_buffer[784] ), .SP(clk_c_enable_659), 
            .CD(n26802), .CK(clk_c), .Q(\data_buffer[792] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i792.GSR = "ENABLED";
    FD1P3IX data_buffer__i788 (.D(\data_buffer[780] ), .SP(clk_c_enable_659), 
            .CD(n26802), .CK(clk_c), .Q(\data_buffer[788] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i788.GSR = "ENABLED";
    FD1P3IX data_buffer__i787 (.D(\data_buffer[779] ), .SP(clk_c_enable_659), 
            .CD(n26803), .CK(clk_c), .Q(\data_buffer[787] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i787.GSR = "ENABLED";
    FD1P3IX data_buffer__i786 (.D(\data_buffer[778] ), .SP(clk_c_enable_659), 
            .CD(n26803), .CK(clk_c), .Q(\data_buffer[786] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i786.GSR = "ENABLED";
    FD1P3IX data_buffer__i785 (.D(\data_buffer[777] ), .SP(clk_c_enable_659), 
            .CD(n26804), .CK(clk_c), .Q(\data_buffer[785] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i785.GSR = "ENABLED";
    FD1P3IX data_buffer__i784 (.D(\data_buffer[776] ), .SP(clk_c_enable_659), 
            .CD(n26803), .CK(clk_c), .Q(\data_buffer[784] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i784.GSR = "ENABLED";
    FD1P3IX data_buffer__i780 (.D(\data_buffer[772] ), .SP(clk_c_enable_659), 
            .CD(n26802), .CK(clk_c), .Q(\data_buffer[780] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i780.GSR = "ENABLED";
    FD1P3IX data_buffer__i779 (.D(\data_buffer[771] ), .SP(clk_c_enable_659), 
            .CD(n26802), .CK(clk_c), .Q(\data_buffer[779] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i779.GSR = "ENABLED";
    FD1P3IX data_buffer__i778 (.D(\data_buffer[770] ), .SP(clk_c_enable_659), 
            .CD(n26799), .CK(clk_c), .Q(\data_buffer[778] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i778.GSR = "ENABLED";
    FD1P3IX data_buffer__i777 (.D(\data_buffer[769] ), .SP(clk_c_enable_659), 
            .CD(n26799), .CK(clk_c), .Q(\data_buffer[777] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i777.GSR = "ENABLED";
    FD1P3IX data_buffer__i776 (.D(\data_buffer[768] ), .SP(clk_c_enable_659), 
            .CD(n26803), .CK(clk_c), .Q(\data_buffer[776] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i776.GSR = "ENABLED";
    FD1P3IX data_buffer__i772 (.D(\data_buffer[764] ), .SP(clk_c_enable_659), 
            .CD(n26804), .CK(clk_c), .Q(\data_buffer[772] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i772.GSR = "ENABLED";
    FD1P3IX data_buffer__i771 (.D(\data_buffer[763] ), .SP(clk_c_enable_659), 
            .CD(n26799), .CK(clk_c), .Q(\data_buffer[771] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i771.GSR = "ENABLED";
    FD1P3IX data_buffer__i770 (.D(\data_buffer[762] ), .SP(clk_c_enable_659), 
            .CD(n26803), .CK(clk_c), .Q(\data_buffer[770] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i770.GSR = "ENABLED";
    FD1P3IX data_buffer__i769 (.D(\data_buffer[761] ), .SP(clk_c_enable_659), 
            .CD(n26804), .CK(clk_c), .Q(\data_buffer[769] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i769.GSR = "ENABLED";
    FD1P3IX data_buffer__i768 (.D(\data_buffer[760] ), .SP(clk_c_enable_659), 
            .CD(n26799), .CK(clk_c), .Q(\data_buffer[768] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i768.GSR = "ENABLED";
    FD1P3IX data_buffer__i764 (.D(\data_buffer[756] ), .SP(clk_c_enable_659), 
            .CD(n26799), .CK(clk_c), .Q(\data_buffer[764] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i764.GSR = "ENABLED";
    FD1P3IX data_buffer__i763 (.D(\data_buffer[755] ), .SP(clk_c_enable_659), 
            .CD(n26799), .CK(clk_c), .Q(\data_buffer[763] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i763.GSR = "ENABLED";
    FD1P3IX data_buffer__i762 (.D(\data_buffer[754] ), .SP(clk_c_enable_659), 
            .CD(n26802), .CK(clk_c), .Q(\data_buffer[762] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i762.GSR = "ENABLED";
    FD1P3IX data_buffer__i761 (.D(\data_buffer[753] ), .SP(clk_c_enable_659), 
            .CD(n26802), .CK(clk_c), .Q(\data_buffer[761] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i761.GSR = "ENABLED";
    FD1P3IX data_buffer__i760 (.D(\data_buffer[752] ), .SP(clk_c_enable_659), 
            .CD(n26804), .CK(clk_c), .Q(\data_buffer[760] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i760.GSR = "ENABLED";
    FD1P3IX data_buffer__i756 (.D(\data_buffer[748] ), .SP(clk_c_enable_659), 
            .CD(n26804), .CK(clk_c), .Q(\data_buffer[756] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i756.GSR = "ENABLED";
    FD1P3IX data_buffer__i755 (.D(\data_buffer[747] ), .SP(clk_c_enable_659), 
            .CD(n26804), .CK(clk_c), .Q(\data_buffer[755] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i755.GSR = "ENABLED";
    FD1P3IX data_buffer__i754 (.D(\data_buffer[746] ), .SP(clk_c_enable_659), 
            .CD(n26804), .CK(clk_c), .Q(\data_buffer[754] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i754.GSR = "ENABLED";
    FD1P3IX data_buffer__i753 (.D(\data_buffer[745] ), .SP(clk_c_enable_659), 
            .CD(n26802), .CK(clk_c), .Q(\data_buffer[753] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i753.GSR = "ENABLED";
    FD1P3IX data_buffer__i752 (.D(\data_buffer[744] ), .SP(clk_c_enable_659), 
            .CD(n26803), .CK(clk_c), .Q(\data_buffer[752] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i752.GSR = "ENABLED";
    FD1P3IX data_buffer__i748 (.D(\data_buffer[740] ), .SP(clk_c_enable_659), 
            .CD(n26804), .CK(clk_c), .Q(\data_buffer[748] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i748.GSR = "ENABLED";
    FD1P3IX data_buffer__i747 (.D(\data_buffer[739] ), .SP(clk_c_enable_659), 
            .CD(n26802), .CK(clk_c), .Q(\data_buffer[747] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i747.GSR = "ENABLED";
    FD1P3IX data_buffer__i746 (.D(\data_buffer[738] ), .SP(clk_c_enable_659), 
            .CD(n26803), .CK(clk_c), .Q(\data_buffer[746] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i746.GSR = "ENABLED";
    FD1P3IX data_buffer__i745 (.D(\data_buffer[737] ), .SP(clk_c_enable_659), 
            .CD(n26805), .CK(clk_c), .Q(\data_buffer[745] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i745.GSR = "ENABLED";
    FD1P3IX data_buffer__i744 (.D(\data_buffer[736] ), .SP(clk_c_enable_659), 
            .CD(n26805), .CK(clk_c), .Q(\data_buffer[744] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i744.GSR = "ENABLED";
    FD1P3IX data_buffer__i740 (.D(\data_buffer[732] ), .SP(clk_c_enable_659), 
            .CD(n26798), .CK(clk_c), .Q(\data_buffer[740] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i740.GSR = "ENABLED";
    FD1P3IX data_buffer__i739 (.D(\data_buffer[731] ), .SP(clk_c_enable_659), 
            .CD(n26799), .CK(clk_c), .Q(\data_buffer[739] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i739.GSR = "ENABLED";
    FD1P3IX data_buffer__i738 (.D(\data_buffer[730] ), .SP(clk_c_enable_659), 
            .CD(n26797), .CK(clk_c), .Q(\data_buffer[738] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i738.GSR = "ENABLED";
    FD1P3IX data_buffer__i737 (.D(\data_buffer[729] ), .SP(clk_c_enable_659), 
            .CD(n26802), .CK(clk_c), .Q(\data_buffer[737] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i737.GSR = "ENABLED";
    FD1P3IX data_buffer__i736 (.D(\data_buffer[728] ), .SP(clk_c_enable_659), 
            .CD(n26805), .CK(clk_c), .Q(\data_buffer[736] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i736.GSR = "ENABLED";
    FD1P3IX data_buffer__i732 (.D(\data_buffer[724] ), .SP(clk_c_enable_659), 
            .CD(n26797), .CK(clk_c), .Q(\data_buffer[732] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i732.GSR = "ENABLED";
    FD1P3IX data_buffer__i731 (.D(\data_buffer[723] ), .SP(clk_c_enable_659), 
            .CD(n26799), .CK(clk_c), .Q(\data_buffer[731] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i731.GSR = "ENABLED";
    FD1P3IX data_buffer__i730 (.D(\data_buffer[722] ), .SP(clk_c_enable_659), 
            .CD(n26794), .CK(clk_c), .Q(\data_buffer[730] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i730.GSR = "ENABLED";
    FD1P3IX data_buffer__i729 (.D(\data_buffer[721] ), .SP(clk_c_enable_659), 
            .CD(n26794), .CK(clk_c), .Q(\data_buffer[729] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i729.GSR = "ENABLED";
    FD1P3IX data_buffer__i728 (.D(\data_buffer[720] ), .SP(clk_c_enable_659), 
            .CD(n26794), .CK(clk_c), .Q(\data_buffer[728] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i728.GSR = "ENABLED";
    FD1P3IX data_buffer__i724 (.D(\data_buffer[716] ), .SP(clk_c_enable_659), 
            .CD(n26794), .CK(clk_c), .Q(\data_buffer[724] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i724.GSR = "ENABLED";
    FD1P3IX data_buffer__i723 (.D(\data_buffer[715] ), .SP(clk_c_enable_659), 
            .CD(n26794), .CK(clk_c), .Q(\data_buffer[723] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i723.GSR = "ENABLED";
    FD1P3IX data_buffer__i722 (.D(\data_buffer[714] ), .SP(clk_c_enable_659), 
            .CD(n26794), .CK(clk_c), .Q(\data_buffer[722] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i722.GSR = "ENABLED";
    FD1P3IX data_buffer__i721 (.D(\data_buffer[713] ), .SP(clk_c_enable_659), 
            .CD(n26794), .CK(clk_c), .Q(\data_buffer[721] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i721.GSR = "ENABLED";
    FD1P3IX data_buffer__i720 (.D(\data_buffer[712] ), .SP(clk_c_enable_659), 
            .CD(n26794), .CK(clk_c), .Q(\data_buffer[720] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i720.GSR = "ENABLED";
    FD1P3IX data_buffer__i716 (.D(\data_buffer[708] ), .SP(clk_c_enable_659), 
            .CD(n26794), .CK(clk_c), .Q(\data_buffer[716] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i716.GSR = "ENABLED";
    FD1P3IX data_buffer__i715 (.D(\data_buffer[707] ), .SP(clk_c_enable_659), 
            .CD(n26794), .CK(clk_c), .Q(\data_buffer[715] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i715.GSR = "ENABLED";
    FD1P3IX data_buffer__i714 (.D(\data_buffer[706] ), .SP(clk_c_enable_659), 
            .CD(n26794), .CK(clk_c), .Q(\data_buffer[714] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i714.GSR = "ENABLED";
    FD1P3IX data_buffer__i713 (.D(\data_buffer[705] ), .SP(clk_c_enable_659), 
            .CD(n26794), .CK(clk_c), .Q(\data_buffer[713] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i713.GSR = "ENABLED";
    FD1P3IX data_buffer__i712 (.D(\data_buffer[704] ), .SP(clk_c_enable_659), 
            .CD(n26799), .CK(clk_c), .Q(\data_buffer[712] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i712.GSR = "ENABLED";
    FD1P3IX data_buffer__i708 (.D(\data_buffer[700] ), .SP(clk_c_enable_659), 
            .CD(n26799), .CK(clk_c), .Q(\data_buffer[708] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i708.GSR = "ENABLED";
    FD1P3IX data_buffer__i707 (.D(\data_buffer[699] ), .SP(clk_c_enable_659), 
            .CD(n26799), .CK(clk_c), .Q(\data_buffer[707] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i707.GSR = "ENABLED";
    FD1P3IX data_buffer__i706 (.D(\data_buffer[698] ), .SP(clk_c_enable_659), 
            .CD(n26799), .CK(clk_c), .Q(\data_buffer[706] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i706.GSR = "ENABLED";
    FD1P3IX data_buffer__i705 (.D(\data_buffer[697] ), .SP(clk_c_enable_659), 
            .CD(n26799), .CK(clk_c), .Q(\data_buffer[705] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i705.GSR = "ENABLED";
    FD1P3IX data_buffer__i704 (.D(\data_buffer[696] ), .SP(clk_c_enable_659), 
            .CD(n26799), .CK(clk_c), .Q(\data_buffer[704] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i704.GSR = "ENABLED";
    FD1P3IX data_buffer__i700 (.D(\data_buffer[692] ), .SP(clk_c_enable_659), 
            .CD(n26799), .CK(clk_c), .Q(\data_buffer[700] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i700.GSR = "ENABLED";
    FD1P3IX data_buffer__i699 (.D(\data_buffer[691] ), .SP(clk_c_enable_659), 
            .CD(n26799), .CK(clk_c), .Q(\data_buffer[699] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i699.GSR = "ENABLED";
    FD1P3IX data_buffer__i698 (.D(\data_buffer[690] ), .SP(clk_c_enable_659), 
            .CD(n26799), .CK(clk_c), .Q(\data_buffer[698] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i698.GSR = "ENABLED";
    FD1P3IX data_buffer__i697 (.D(\data_buffer[689] ), .SP(clk_c_enable_659), 
            .CD(n26799), .CK(clk_c), .Q(\data_buffer[697] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i697.GSR = "ENABLED";
    FD1P3IX data_buffer__i696 (.D(\data_buffer[688] ), .SP(clk_c_enable_659), 
            .CD(n26794), .CK(clk_c), .Q(\data_buffer[696] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i696.GSR = "ENABLED";
    FD1P3IX data_buffer__i692 (.D(\data_buffer[684] ), .SP(clk_c_enable_659), 
            .CD(n26799), .CK(clk_c), .Q(\data_buffer[692] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i692.GSR = "ENABLED";
    FD1P3IX data_buffer__i691 (.D(\data_buffer[683] ), .SP(clk_c_enable_659), 
            .CD(n26794), .CK(clk_c), .Q(\data_buffer[691] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i691.GSR = "ENABLED";
    FD1P3IX data_buffer__i690 (.D(\data_buffer[682] ), .SP(clk_c_enable_659), 
            .CD(n26794), .CK(clk_c), .Q(\data_buffer[690] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i690.GSR = "ENABLED";
    FD1P3IX data_buffer__i689 (.D(\data_buffer[681] ), .SP(clk_c_enable_659), 
            .CD(n26799), .CK(clk_c), .Q(\data_buffer[689] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i689.GSR = "ENABLED";
    FD1P3IX data_buffer__i688 (.D(\data_buffer[680] ), .SP(clk_c_enable_659), 
            .CD(n26794), .CK(clk_c), .Q(\data_buffer[688] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i688.GSR = "ENABLED";
    FD1P3IX data_buffer__i684 (.D(\data_buffer[676] ), .SP(clk_c_enable_659), 
            .CD(n26794), .CK(clk_c), .Q(\data_buffer[684] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i684.GSR = "ENABLED";
    FD1P3IX data_buffer__i683 (.D(\data_buffer[675] ), .SP(clk_c_enable_659), 
            .CD(n26799), .CK(clk_c), .Q(\data_buffer[683] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i683.GSR = "ENABLED";
    FD1P3IX data_buffer__i682 (.D(\data_buffer[674] ), .SP(clk_c_enable_659), 
            .CD(n26794), .CK(clk_c), .Q(\data_buffer[682] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i682.GSR = "ENABLED";
    FD1P3IX data_buffer__i681 (.D(\data_buffer[673] ), .SP(clk_c_enable_659), 
            .CD(n26799), .CK(clk_c), .Q(\data_buffer[681] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i681.GSR = "ENABLED";
    FD1P3IX data_buffer__i680 (.D(\data_buffer[672] ), .SP(clk_c_enable_659), 
            .CD(n26794), .CK(clk_c), .Q(\data_buffer[680] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i680.GSR = "ENABLED";
    FD1P3IX data_buffer__i676 (.D(\data_buffer[668] ), .SP(clk_c_enable_659), 
            .CD(n26794), .CK(clk_c), .Q(\data_buffer[676] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i676.GSR = "ENABLED";
    FD1P3IX data_buffer__i675 (.D(\data_buffer[667] ), .SP(clk_c_enable_659), 
            .CD(n26799), .CK(clk_c), .Q(\data_buffer[675] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i675.GSR = "ENABLED";
    FD1P3IX data_buffer__i674 (.D(\data_buffer[666] ), .SP(clk_c_enable_659), 
            .CD(n26794), .CK(clk_c), .Q(\data_buffer[674] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i674.GSR = "ENABLED";
    FD1P3IX data_buffer__i673 (.D(\data_buffer[665] ), .SP(clk_c_enable_659), 
            .CD(n26799), .CK(clk_c), .Q(\data_buffer[673] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i673.GSR = "ENABLED";
    FD1P3IX data_buffer__i672 (.D(\data_buffer[664] ), .SP(clk_c_enable_659), 
            .CD(n26794), .CK(clk_c), .Q(\data_buffer[672] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i672.GSR = "ENABLED";
    FD1P3IX data_buffer__i668 (.D(\data_buffer[660] ), .SP(clk_c_enable_659), 
            .CD(n26799), .CK(clk_c), .Q(\data_buffer[668] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i668.GSR = "ENABLED";
    FD1P3IX data_buffer__i667 (.D(\data_buffer[659] ), .SP(clk_c_enable_659), 
            .CD(n26805), .CK(clk_c), .Q(\data_buffer[667] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i667.GSR = "ENABLED";
    FD1P3IX data_buffer__i666 (.D(\data_buffer[658] ), .SP(clk_c_enable_659), 
            .CD(n26805), .CK(clk_c), .Q(\data_buffer[666] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i666.GSR = "ENABLED";
    FD1P3IX data_buffer__i665 (.D(\data_buffer[657] ), .SP(clk_c_enable_659), 
            .CD(n26803), .CK(clk_c), .Q(\data_buffer[665] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i665.GSR = "ENABLED";
    FD1P3IX data_buffer__i664 (.D(\data_buffer[656] ), .SP(clk_c_enable_659), 
            .CD(n26805), .CK(clk_c), .Q(\data_buffer[664] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i664.GSR = "ENABLED";
    FD1P3IX data_buffer__i660 (.D(\data_buffer[652] ), .SP(clk_c_enable_659), 
            .CD(n26799), .CK(clk_c), .Q(\data_buffer[660] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i660.GSR = "ENABLED";
    FD1P3IX data_buffer__i659 (.D(\data_buffer[651] ), .SP(clk_c_enable_659), 
            .CD(n26801), .CK(clk_c), .Q(\data_buffer[659] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i659.GSR = "ENABLED";
    FD1P3IX data_buffer__i658 (.D(\data_buffer[650] ), .SP(clk_c_enable_659), 
            .CD(n26801), .CK(clk_c), .Q(\data_buffer[658] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i658.GSR = "ENABLED";
    FD1P3IX data_buffer__i657 (.D(\data_buffer[649] ), .SP(clk_c_enable_659), 
            .CD(n26799), .CK(clk_c), .Q(\data_buffer[657] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i657.GSR = "ENABLED";
    FD1P3IX data_buffer__i656 (.D(\data_buffer[648] ), .SP(clk_c_enable_659), 
            .CD(n26799), .CK(clk_c), .Q(\data_buffer[656] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i656.GSR = "ENABLED";
    FD1P3IX data_buffer__i652 (.D(\data_buffer[644] ), .SP(clk_c_enable_659), 
            .CD(n26801), .CK(clk_c), .Q(\data_buffer[652] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i652.GSR = "ENABLED";
    FD1P3IX data_buffer__i651 (.D(\data_buffer[643] ), .SP(clk_c_enable_659), 
            .CD(n26801), .CK(clk_c), .Q(\data_buffer[651] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i651.GSR = "ENABLED";
    FD1P3IX data_buffer__i650 (.D(\data_buffer[642] ), .SP(clk_c_enable_659), 
            .CD(n26801), .CK(clk_c), .Q(\data_buffer[650] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i650.GSR = "ENABLED";
    FD1P3IX data_buffer__i649 (.D(\data_buffer[641] ), .SP(clk_c_enable_659), 
            .CD(n26801), .CK(clk_c), .Q(\data_buffer[649] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i649.GSR = "ENABLED";
    FD1P3IX data_buffer__i648 (.D(\data_buffer[640] ), .SP(clk_c_enable_659), 
            .CD(n26801), .CK(clk_c), .Q(\data_buffer[648] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i648.GSR = "ENABLED";
    FD1P3IX data_buffer__i644 (.D(\data_buffer[636] ), .SP(clk_c_enable_659), 
            .CD(n26801), .CK(clk_c), .Q(\data_buffer[644] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i644.GSR = "ENABLED";
    FD1P3IX data_buffer__i643 (.D(\data_buffer[635] ), .SP(clk_c_enable_659), 
            .CD(n26801), .CK(clk_c), .Q(\data_buffer[643] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i643.GSR = "ENABLED";
    FD1P3IX data_buffer__i642 (.D(\data_buffer[634] ), .SP(clk_c_enable_659), 
            .CD(n26801), .CK(clk_c), .Q(\data_buffer[642] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i642.GSR = "ENABLED";
    FD1P3IX data_buffer__i641 (.D(\data_buffer[633] ), .SP(clk_c_enable_659), 
            .CD(n26801), .CK(clk_c), .Q(\data_buffer[641] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i641.GSR = "ENABLED";
    FD1P3IX data_buffer__i640 (.D(\data_buffer[632] ), .SP(clk_c_enable_659), 
            .CD(n26801), .CK(clk_c), .Q(\data_buffer[640] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i640.GSR = "ENABLED";
    FD1P3IX data_buffer__i636 (.D(\data_buffer[628] ), .SP(clk_c_enable_659), 
            .CD(n26801), .CK(clk_c), .Q(\data_buffer[636] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i636.GSR = "ENABLED";
    FD1P3IX data_buffer__i635 (.D(\data_buffer[627] ), .SP(clk_c_enable_659), 
            .CD(n26803), .CK(clk_c), .Q(\data_buffer[635] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i635.GSR = "ENABLED";
    FD1P3IX data_buffer__i634 (.D(\data_buffer[626] ), .SP(clk_c_enable_659), 
            .CD(n26803), .CK(clk_c), .Q(\data_buffer[634] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i634.GSR = "ENABLED";
    FD1P3IX data_buffer__i633 (.D(\data_buffer[625] ), .SP(clk_c_enable_659), 
            .CD(n26803), .CK(clk_c), .Q(\data_buffer[633] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i633.GSR = "ENABLED";
    FD1P3IX data_buffer__i632 (.D(\data_buffer[624] ), .SP(clk_c_enable_659), 
            .CD(n26805), .CK(clk_c), .Q(\data_buffer[632] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i632.GSR = "ENABLED";
    FD1P3IX data_buffer__i628 (.D(\data_buffer[620] ), .SP(clk_c_enable_659), 
            .CD(n26797), .CK(clk_c), .Q(\data_buffer[628] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i628.GSR = "ENABLED";
    FD1P3IX data_buffer__i627 (.D(\data_buffer[619] ), .SP(clk_c_enable_659), 
            .CD(n26800), .CK(clk_c), .Q(\data_buffer[627] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i627.GSR = "ENABLED";
    FD1P3IX data_buffer__i626 (.D(\data_buffer[618] ), .SP(clk_c_enable_659), 
            .CD(n26800), .CK(clk_c), .Q(\data_buffer[626] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i626.GSR = "ENABLED";
    FD1P3IX data_buffer__i625 (.D(\data_buffer[617] ), .SP(clk_c_enable_659), 
            .CD(n26800), .CK(clk_c), .Q(\data_buffer[625] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i625.GSR = "ENABLED";
    FD1P3IX data_buffer__i624 (.D(\data_buffer[616] ), .SP(clk_c_enable_659), 
            .CD(n26800), .CK(clk_c), .Q(\data_buffer[624] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i624.GSR = "ENABLED";
    FD1P3IX data_buffer__i620 (.D(\data_buffer[612] ), .SP(clk_c_enable_659), 
            .CD(n26800), .CK(clk_c), .Q(\data_buffer[620] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i620.GSR = "ENABLED";
    FD1P3IX data_buffer__i619 (.D(\data_buffer[611] ), .SP(clk_c_enable_659), 
            .CD(n26799), .CK(clk_c), .Q(\data_buffer[619] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i619.GSR = "ENABLED";
    FD1P3IX data_buffer__i618 (.D(\data_buffer[610] ), .SP(clk_c_enable_659), 
            .CD(n26802), .CK(clk_c), .Q(\data_buffer[618] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i618.GSR = "ENABLED";
    FD1P3IX data_buffer__i617 (.D(\data_buffer[609] ), .SP(clk_c_enable_659), 
            .CD(n26797), .CK(clk_c), .Q(\data_buffer[617] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i617.GSR = "ENABLED";
    FD1P3IX data_buffer__i616 (.D(\data_buffer[608] ), .SP(clk_c_enable_659), 
            .CD(n26802), .CK(clk_c), .Q(\data_buffer[616] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i616.GSR = "ENABLED";
    FD1P3IX data_buffer__i612 (.D(\data_buffer[604] ), .SP(clk_c_enable_659), 
            .CD(n26798), .CK(clk_c), .Q(\data_buffer[612] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i612.GSR = "ENABLED";
    FD1P3IX data_buffer__i611 (.D(\data_buffer[603] ), .SP(clk_c_enable_659), 
            .CD(n26805), .CK(clk_c), .Q(\data_buffer[611] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i611.GSR = "ENABLED";
    FD1P3IX data_buffer__i610 (.D(\data_buffer[602] ), .SP(clk_c_enable_659), 
            .CD(n26799), .CK(clk_c), .Q(\data_buffer[610] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i610.GSR = "ENABLED";
    FD1P3IX data_buffer__i609 (.D(\data_buffer[601] ), .SP(clk_c_enable_659), 
            .CD(n26798), .CK(clk_c), .Q(\data_buffer[609] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i609.GSR = "ENABLED";
    FD1P3IX data_buffer__i608 (.D(\data_buffer[600] ), .SP(clk_c_enable_659), 
            .CD(n26798), .CK(clk_c), .Q(\data_buffer[608] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i608.GSR = "ENABLED";
    FD1P3IX data_buffer__i604 (.D(\data_buffer[596] ), .SP(clk_c_enable_659), 
            .CD(n26805), .CK(clk_c), .Q(\data_buffer[604] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i604.GSR = "ENABLED";
    FD1P3IX data_buffer__i603 (.D(\data_buffer[595] ), .SP(clk_c_enable_659), 
            .CD(n26798), .CK(clk_c), .Q(\data_buffer[603] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i603.GSR = "ENABLED";
    FD1P3IX data_buffer__i602 (.D(\data_buffer[594] ), .SP(clk_c_enable_659), 
            .CD(n26805), .CK(clk_c), .Q(\data_buffer[602] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i602.GSR = "ENABLED";
    FD1P3IX data_buffer__i601 (.D(\data_buffer[593] ), .SP(clk_c_enable_659), 
            .CD(n26803), .CK(clk_c), .Q(\data_buffer[601] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i601.GSR = "ENABLED";
    FD1P3IX data_buffer__i600 (.D(\data_buffer[592] ), .SP(clk_c_enable_659), 
            .CD(n26805), .CK(clk_c), .Q(\data_buffer[600] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i600.GSR = "ENABLED";
    FD1P3IX data_buffer__i596 (.D(\data_buffer[588] ), .SP(clk_c_enable_659), 
            .CD(n26803), .CK(clk_c), .Q(\data_buffer[596] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i596.GSR = "ENABLED";
    FD1P3IX data_buffer__i595 (.D(\data_buffer[587] ), .SP(clk_c_enable_659), 
            .CD(n26805), .CK(clk_c), .Q(\data_buffer[595] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i595.GSR = "ENABLED";
    FD1P3IX data_buffer__i594 (.D(\data_buffer[586] ), .SP(clk_c_enable_659), 
            .CD(n26803), .CK(clk_c), .Q(\data_buffer[594] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i594.GSR = "ENABLED";
    FD1P3IX data_buffer__i593 (.D(\data_buffer[585] ), .SP(clk_c_enable_659), 
            .CD(n26805), .CK(clk_c), .Q(\data_buffer[593] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i593.GSR = "ENABLED";
    FD1P3IX data_buffer__i592 (.D(\data_buffer[584] ), .SP(clk_c_enable_659), 
            .CD(n26803), .CK(clk_c), .Q(\data_buffer[592] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i592.GSR = "ENABLED";
    FD1P3IX data_buffer__i588 (.D(\data_buffer[580] ), .SP(clk_c_enable_659), 
            .CD(n26805), .CK(clk_c), .Q(\data_buffer[588] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i588.GSR = "ENABLED";
    FD1P3IX data_buffer__i587 (.D(\data_buffer[579] ), .SP(clk_c_enable_659), 
            .CD(n26805), .CK(clk_c), .Q(\data_buffer[587] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i587.GSR = "ENABLED";
    FD1P3IX data_buffer__i586 (.D(\data_buffer[578] ), .SP(clk_c_enable_659), 
            .CD(n26797), .CK(clk_c), .Q(\data_buffer[586] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i586.GSR = "ENABLED";
    FD1P3IX data_buffer__i585 (.D(\data_buffer[577] ), .SP(clk_c_enable_659), 
            .CD(n26805), .CK(clk_c), .Q(\data_buffer[585] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i585.GSR = "ENABLED";
    FD1P3IX data_buffer__i584 (.D(\data_buffer[576] ), .SP(clk_c_enable_659), 
            .CD(n26805), .CK(clk_c), .Q(\data_buffer[584] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i584.GSR = "ENABLED";
    FD1P3IX data_buffer__i580 (.D(\data_buffer[572] ), .SP(clk_c_enable_659), 
            .CD(n26805), .CK(clk_c), .Q(\data_buffer[580] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i580.GSR = "ENABLED";
    FD1P3IX data_buffer__i579 (.D(\data_buffer[571] ), .SP(clk_c_enable_659), 
            .CD(n26797), .CK(clk_c), .Q(\data_buffer[579] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i579.GSR = "ENABLED";
    FD1P3IX data_buffer__i578 (.D(\data_buffer[570] ), .SP(clk_c_enable_659), 
            .CD(n26801), .CK(clk_c), .Q(\data_buffer[578] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i578.GSR = "ENABLED";
    FD1P3IX data_buffer__i577 (.D(\data_buffer[569] ), .SP(clk_c_enable_659), 
            .CD(n26805), .CK(clk_c), .Q(\data_buffer[577] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i577.GSR = "ENABLED";
    FD1P3IX data_buffer__i576 (.D(\data_buffer[568] ), .SP(clk_c_enable_659), 
            .CD(n26801), .CK(clk_c), .Q(\data_buffer[576] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i576.GSR = "ENABLED";
    FD1P3IX data_buffer__i572 (.D(\data_buffer[564] ), .SP(clk_c_enable_659), 
            .CD(n26801), .CK(clk_c), .Q(\data_buffer[572] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i572.GSR = "ENABLED";
    FD1P3IX data_buffer__i571 (.D(\data_buffer[563] ), .SP(clk_c_enable_659), 
            .CD(n26805), .CK(clk_c), .Q(\data_buffer[571] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i571.GSR = "ENABLED";
    FD1P3IX data_buffer__i570 (.D(\data_buffer[562] ), .SP(clk_c_enable_659), 
            .CD(n26801), .CK(clk_c), .Q(\data_buffer[570] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i570.GSR = "ENABLED";
    FD1P3IX data_buffer__i569 (.D(\data_buffer[561] ), .SP(clk_c_enable_659), 
            .CD(n26801), .CK(clk_c), .Q(\data_buffer[569] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i569.GSR = "ENABLED";
    FD1P3IX data_buffer__i568 (.D(\data_buffer[560] ), .SP(clk_c_enable_659), 
            .CD(n26805), .CK(clk_c), .Q(\data_buffer[568] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i568.GSR = "ENABLED";
    FD1P3IX data_buffer__i564 (.D(\data_buffer[556] ), .SP(clk_c_enable_659), 
            .CD(n26799), .CK(clk_c), .Q(\data_buffer[564] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i564.GSR = "ENABLED";
    FD1P3IX data_buffer__i563 (.D(\data_buffer[555] ), .SP(clk_c_enable_659), 
            .CD(n26799), .CK(clk_c), .Q(\data_buffer[563] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i563.GSR = "ENABLED";
    FD1P3IX data_buffer__i562 (.D(\data_buffer[554] ), .SP(clk_c_enable_659), 
            .CD(n26802), .CK(clk_c), .Q(\data_buffer[562] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i562.GSR = "ENABLED";
    FD1P3IX data_buffer__i561 (.D(\data_buffer[553] ), .SP(clk_c_enable_659), 
            .CD(n26805), .CK(clk_c), .Q(\data_buffer[561] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i561.GSR = "ENABLED";
    FD1P3IX data_buffer__i560 (.D(\data_buffer[552] ), .SP(clk_c_enable_659), 
            .CD(n26799), .CK(clk_c), .Q(\data_buffer[560] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i560.GSR = "ENABLED";
    FD1P3IX data_buffer__i556 (.D(\data_buffer[548] ), .SP(clk_c_enable_659), 
            .CD(n26801), .CK(clk_c), .Q(\data_buffer[556] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i556.GSR = "ENABLED";
    FD1P3IX data_buffer__i555 (.D(\data_buffer[547] ), .SP(clk_c_enable_659), 
            .CD(n26805), .CK(clk_c), .Q(\data_buffer[555] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i555.GSR = "ENABLED";
    FD1P3IX data_buffer__i554 (.D(\data_buffer[546] ), .SP(clk_c_enable_659), 
            .CD(n26801), .CK(clk_c), .Q(\data_buffer[554] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i554.GSR = "ENABLED";
    FD1P3IX data_buffer__i553 (.D(\data_buffer[545] ), .SP(clk_c_enable_659), 
            .CD(n26802), .CK(clk_c), .Q(\data_buffer[553] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i553.GSR = "ENABLED";
    FD1P3IX data_buffer__i552 (.D(\data_buffer[544] ), .SP(clk_c_enable_659), 
            .CD(n26798), .CK(clk_c), .Q(\data_buffer[552] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i552.GSR = "ENABLED";
    FD1P3IX data_buffer__i548 (.D(\data_buffer[540] ), .SP(clk_c_enable_659), 
            .CD(n26794), .CK(clk_c), .Q(\data_buffer[548] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i548.GSR = "ENABLED";
    FD1P3IX data_buffer__i547 (.D(\data_buffer[539] ), .SP(clk_c_enable_659), 
            .CD(n26794), .CK(clk_c), .Q(\data_buffer[547] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i547.GSR = "ENABLED";
    FD1P3IX data_buffer__i546 (.D(\data_buffer[538] ), .SP(clk_c_enable_659), 
            .CD(n26794), .CK(clk_c), .Q(\data_buffer[546] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i546.GSR = "ENABLED";
    FD1P3IX data_buffer__i545 (.D(\data_buffer[537] ), .SP(clk_c_enable_659), 
            .CD(n26794), .CK(clk_c), .Q(\data_buffer[545] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i545.GSR = "ENABLED";
    FD1P3IX data_buffer__i544 (.D(\data_buffer[536] ), .SP(clk_c_enable_659), 
            .CD(n26794), .CK(clk_c), .Q(\data_buffer[544] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i544.GSR = "ENABLED";
    FD1P3IX data_buffer__i540 (.D(\data_buffer[532] ), .SP(clk_c_enable_659), 
            .CD(n26794), .CK(clk_c), .Q(\data_buffer[540] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i540.GSR = "ENABLED";
    FD1P3IX data_buffer__i539 (.D(\data_buffer[531] ), .SP(clk_c_enable_659), 
            .CD(n26802), .CK(clk_c), .Q(\data_buffer[539] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i539.GSR = "ENABLED";
    FD1P3IX data_buffer__i538 (.D(\data_buffer[530] ), .SP(clk_c_enable_659), 
            .CD(n26794), .CK(clk_c), .Q(\data_buffer[538] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i538.GSR = "ENABLED";
    FD1P3IX data_buffer__i537 (.D(\data_buffer[529] ), .SP(clk_c_enable_659), 
            .CD(n26802), .CK(clk_c), .Q(\data_buffer[537] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i537.GSR = "ENABLED";
    FD1P3IX data_buffer__i536 (.D(\data_buffer[528] ), .SP(clk_c_enable_659), 
            .CD(n26799), .CK(clk_c), .Q(\data_buffer[536] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i536.GSR = "ENABLED";
    FD1P3IX data_buffer__i532 (.D(\data_buffer[524] ), .SP(clk_c_enable_659), 
            .CD(n26799), .CK(clk_c), .Q(\data_buffer[532] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i532.GSR = "ENABLED";
    FD1P3IX data_buffer__i531 (.D(\data_buffer[523] ), .SP(clk_c_enable_659), 
            .CD(n26803), .CK(clk_c), .Q(\data_buffer[531] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i531.GSR = "ENABLED";
    FD1P3IX data_buffer__i530 (.D(\data_buffer[522] ), .SP(clk_c_enable_659), 
            .CD(n26799), .CK(clk_c), .Q(\data_buffer[530] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i530.GSR = "ENABLED";
    FD1P3IX data_buffer__i529 (.D(\data_buffer[521] ), .SP(clk_c_enable_659), 
            .CD(n26799), .CK(clk_c), .Q(\data_buffer[529] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i529.GSR = "ENABLED";
    FD1P3IX data_buffer__i528 (.D(\data_buffer[520] ), .SP(clk_c_enable_659), 
            .CD(n26794), .CK(clk_c), .Q(\data_buffer[528] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i528.GSR = "ENABLED";
    FD1P3IX data_buffer__i524 (.D(\data_buffer[516] ), .SP(clk_c_enable_659), 
            .CD(n26805), .CK(clk_c), .Q(\data_buffer[524] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i524.GSR = "ENABLED";
    FD1P3IX data_buffer__i523 (.D(\data_buffer[515] ), .SP(clk_c_enable_659), 
            .CD(n26802), .CK(clk_c), .Q(\data_buffer[523] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i523.GSR = "ENABLED";
    FD1P3IX data_buffer__i522 (.D(\data_buffer[514] ), .SP(clk_c_enable_659), 
            .CD(n26802), .CK(clk_c), .Q(\data_buffer[522] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i522.GSR = "ENABLED";
    FD1P3IX data_buffer__i521 (.D(\data_buffer[513] ), .SP(clk_c_enable_659), 
            .CD(n26802), .CK(clk_c), .Q(\data_buffer[521] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i521.GSR = "ENABLED";
    FD1P3IX data_buffer__i520 (.D(\data_buffer[512] ), .SP(clk_c_enable_659), 
            .CD(n26799), .CK(clk_c), .Q(\data_buffer[520] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i520.GSR = "ENABLED";
    FD1P3IX data_buffer__i516 (.D(\data_buffer[508] ), .SP(clk_c_enable_659), 
            .CD(n26794), .CK(clk_c), .Q(\data_buffer[516] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i516.GSR = "ENABLED";
    FD1P3IX data_buffer__i515 (.D(\data_buffer[507] ), .SP(clk_c_enable_659), 
            .CD(n26794), .CK(clk_c), .Q(\data_buffer[515] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i515.GSR = "ENABLED";
    FD1P3IX data_buffer__i514 (.D(\data_buffer[506] ), .SP(clk_c_enable_659), 
            .CD(n26794), .CK(clk_c), .Q(\data_buffer[514] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i514.GSR = "ENABLED";
    FD1P3IX data_buffer__i513 (.D(\data_buffer[505] ), .SP(clk_c_enable_659), 
            .CD(n26794), .CK(clk_c), .Q(\data_buffer[513] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i513.GSR = "ENABLED";
    FD1P3IX data_buffer__i512 (.D(\data_buffer[504] ), .SP(clk_c_enable_659), 
            .CD(n26794), .CK(clk_c), .Q(\data_buffer[512] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i512.GSR = "ENABLED";
    FD1P3IX data_buffer__i508 (.D(\data_buffer[500] ), .SP(clk_c_enable_659), 
            .CD(n26794), .CK(clk_c), .Q(\data_buffer[508] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i508.GSR = "ENABLED";
    FD1P3IX data_buffer__i507 (.D(\data_buffer[499] ), .SP(clk_c_enable_659), 
            .CD(n26794), .CK(clk_c), .Q(\data_buffer[507] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i507.GSR = "ENABLED";
    FD1P3IX data_buffer__i506 (.D(\data_buffer[498] ), .SP(clk_c_enable_659), 
            .CD(n26794), .CK(clk_c), .Q(\data_buffer[506] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i506.GSR = "ENABLED";
    FD1P3IX data_buffer__i505 (.D(\data_buffer[497] ), .SP(clk_c_enable_659), 
            .CD(n26794), .CK(clk_c), .Q(\data_buffer[505] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i505.GSR = "ENABLED";
    FD1P3IX data_buffer__i504 (.D(\data_buffer[496] ), .SP(clk_c_enable_659), 
            .CD(n26794), .CK(clk_c), .Q(\data_buffer[504] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i504.GSR = "ENABLED";
    FD1P3IX data_buffer__i500 (.D(\data_buffer[492] ), .SP(clk_c_enable_659), 
            .CD(n26794), .CK(clk_c), .Q(\data_buffer[500] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i500.GSR = "ENABLED";
    FD1P3IX data_buffer__i499 (.D(\data_buffer[491] ), .SP(clk_c_enable_659), 
            .CD(n26799), .CK(clk_c), .Q(\data_buffer[499] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i499.GSR = "ENABLED";
    FD1P3IX data_buffer__i498 (.D(\data_buffer[490] ), .SP(clk_c_enable_659), 
            .CD(n26794), .CK(clk_c), .Q(\data_buffer[498] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i498.GSR = "ENABLED";
    FD1P3IX data_buffer__i497 (.D(\data_buffer[489] ), .SP(clk_c_enable_659), 
            .CD(n26794), .CK(clk_c), .Q(\data_buffer[497] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i497.GSR = "ENABLED";
    FD1P3IX data_buffer__i496 (.D(\data_buffer[488] ), .SP(clk_c_enable_659), 
            .CD(n26794), .CK(clk_c), .Q(\data_buffer[496] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i496.GSR = "ENABLED";
    FD1P3IX data_buffer__i492 (.D(\data_buffer[484] ), .SP(clk_c_enable_659), 
            .CD(n26799), .CK(clk_c), .Q(\data_buffer[492] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i492.GSR = "ENABLED";
    FD1P3IX data_buffer__i491 (.D(\data_buffer[483] ), .SP(clk_c_enable_659), 
            .CD(n26794), .CK(clk_c), .Q(\data_buffer[491] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i491.GSR = "ENABLED";
    FD1P3IX data_buffer__i490 (.D(\data_buffer[482] ), .SP(clk_c_enable_659), 
            .CD(n26795), .CK(clk_c), .Q(\data_buffer[490] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i490.GSR = "ENABLED";
    FD1P3IX data_buffer__i489 (.D(\data_buffer[481] ), .SP(clk_c_enable_659), 
            .CD(n26795), .CK(clk_c), .Q(\data_buffer[489] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i489.GSR = "ENABLED";
    FD1P3IX data_buffer__i488 (.D(\data_buffer[480] ), .SP(clk_c_enable_659), 
            .CD(n26795), .CK(clk_c), .Q(\data_buffer[488] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i488.GSR = "ENABLED";
    FD1P3IX data_buffer__i484 (.D(\data_buffer[476] ), .SP(clk_c_enable_659), 
            .CD(n26795), .CK(clk_c), .Q(\data_buffer[484] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i484.GSR = "ENABLED";
    FD1P3IX data_buffer__i483 (.D(\data_buffer[475] ), .SP(clk_c_enable_659), 
            .CD(n26795), .CK(clk_c), .Q(\data_buffer[483] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i483.GSR = "ENABLED";
    FD1P3IX data_buffer__i482 (.D(\data_buffer[474] ), .SP(clk_c_enable_659), 
            .CD(n26794), .CK(clk_c), .Q(\data_buffer[482] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i482.GSR = "ENABLED";
    FD1P3IX data_buffer__i481 (.D(\data_buffer[473] ), .SP(clk_c_enable_659), 
            .CD(n26795), .CK(clk_c), .Q(\data_buffer[481] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i481.GSR = "ENABLED";
    FD1P3IX data_buffer__i480 (.D(\data_buffer[472] ), .SP(clk_c_enable_659), 
            .CD(n26794), .CK(clk_c), .Q(\data_buffer[480] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i480.GSR = "ENABLED";
    FD1P3IX data_buffer__i476 (.D(\data_buffer[468] ), .SP(clk_c_enable_659), 
            .CD(n26794), .CK(clk_c), .Q(\data_buffer[476] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i476.GSR = "ENABLED";
    FD1P3IX data_buffer__i475 (.D(\data_buffer[467] ), .SP(clk_c_enable_659), 
            .CD(n26795), .CK(clk_c), .Q(\data_buffer[475] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i475.GSR = "ENABLED";
    FD1P3IX data_buffer__i474 (.D(\data_buffer[466] ), .SP(clk_c_enable_659), 
            .CD(n26795), .CK(clk_c), .Q(\data_buffer[474] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i474.GSR = "ENABLED";
    FD1P3IX data_buffer__i473 (.D(\data_buffer[465] ), .SP(clk_c_enable_659), 
            .CD(n26795), .CK(clk_c), .Q(\data_buffer[473] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i473.GSR = "ENABLED";
    FD1P3IX data_buffer__i472 (.D(\data_buffer[464] ), .SP(clk_c_enable_659), 
            .CD(n26795), .CK(clk_c), .Q(\data_buffer[472] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i472.GSR = "ENABLED";
    FD1P3IX data_buffer__i468 (.D(\data_buffer[460] ), .SP(clk_c_enable_659), 
            .CD(n26795), .CK(clk_c), .Q(\data_buffer[468] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i468.GSR = "ENABLED";
    FD1P3IX data_buffer__i467 (.D(\data_buffer[459] ), .SP(clk_c_enable_659), 
            .CD(n26795), .CK(clk_c), .Q(\data_buffer[467] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i467.GSR = "ENABLED";
    FD1P3IX data_buffer__i466 (.D(\data_buffer[458] ), .SP(clk_c_enable_659), 
            .CD(n26795), .CK(clk_c), .Q(\data_buffer[466] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i466.GSR = "ENABLED";
    FD1P3IX data_buffer__i465 (.D(\data_buffer[457] ), .SP(clk_c_enable_659), 
            .CD(n26795), .CK(clk_c), .Q(\data_buffer[465] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i465.GSR = "ENABLED";
    FD1P3IX data_buffer__i464 (.D(\data_buffer[456] ), .SP(clk_c_enable_659), 
            .CD(n26795), .CK(clk_c), .Q(\data_buffer[464] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i464.GSR = "ENABLED";
    FD1P3IX data_buffer__i460 (.D(\data_buffer[452] ), .SP(clk_c_enable_659), 
            .CD(n26795), .CK(clk_c), .Q(\data_buffer[460] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i460.GSR = "ENABLED";
    FD1P3IX data_buffer__i459 (.D(\data_buffer[451] ), .SP(clk_c_enable_659), 
            .CD(n26795), .CK(clk_c), .Q(\data_buffer[459] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i459.GSR = "ENABLED";
    FD1P3IX data_buffer__i458 (.D(\data_buffer[450] ), .SP(clk_c_enable_659), 
            .CD(n26795), .CK(clk_c), .Q(\data_buffer[458] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i458.GSR = "ENABLED";
    FD1P3IX data_buffer__i457 (.D(\data_buffer[449] ), .SP(clk_c_enable_659), 
            .CD(n26795), .CK(clk_c), .Q(\data_buffer[457] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i457.GSR = "ENABLED";
    FD1P3IX data_buffer__i456 (.D(\data_buffer[448] ), .SP(clk_c_enable_659), 
            .CD(n26795), .CK(clk_c), .Q(\data_buffer[456] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i456.GSR = "ENABLED";
    FD1P3IX data_buffer__i452 (.D(\data_buffer[444] ), .SP(clk_c_enable_659), 
            .CD(n26795), .CK(clk_c), .Q(\data_buffer[452] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i452.GSR = "ENABLED";
    FD1P3IX data_buffer__i451 (.D(\data_buffer[443] ), .SP(clk_c_enable_659), 
            .CD(n26795), .CK(clk_c), .Q(\data_buffer[451] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i451.GSR = "ENABLED";
    FD1P3IX data_buffer__i450 (.D(\data_buffer[442] ), .SP(clk_c_enable_659), 
            .CD(n26795), .CK(clk_c), .Q(\data_buffer[450] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i450.GSR = "ENABLED";
    FD1P3IX data_buffer__i449 (.D(\data_buffer[441] ), .SP(clk_c_enable_659), 
            .CD(n26795), .CK(clk_c), .Q(\data_buffer[449] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i449.GSR = "ENABLED";
    FD1P3IX data_buffer__i448 (.D(\data_buffer[440] ), .SP(clk_c_enable_659), 
            .CD(n26795), .CK(clk_c), .Q(\data_buffer[448] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i448.GSR = "ENABLED";
    FD1P3IX data_buffer__i444 (.D(\data_buffer[436] ), .SP(clk_c_enable_659), 
            .CD(n26795), .CK(clk_c), .Q(\data_buffer[444] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i444.GSR = "ENABLED";
    FD1P3IX data_buffer__i443 (.D(\data_buffer[435] ), .SP(clk_c_enable_659), 
            .CD(n26795), .CK(clk_c), .Q(\data_buffer[443] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i443.GSR = "ENABLED";
    FD1P3IX data_buffer__i442 (.D(\data_buffer[434] ), .SP(clk_c_enable_659), 
            .CD(n26795), .CK(clk_c), .Q(\data_buffer[442] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i442.GSR = "ENABLED";
    FD1P3IX data_buffer__i441 (.D(\data_buffer[433] ), .SP(clk_c_enable_659), 
            .CD(n26795), .CK(clk_c), .Q(\data_buffer[441] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i441.GSR = "ENABLED";
    FD1P3IX data_buffer__i440 (.D(\data_buffer[432] ), .SP(clk_c_enable_659), 
            .CD(n26795), .CK(clk_c), .Q(\data_buffer[440] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i440.GSR = "ENABLED";
    FD1P3IX data_buffer__i436 (.D(\data_buffer[428] ), .SP(clk_c_enable_659), 
            .CD(n26795), .CK(clk_c), .Q(\data_buffer[436] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i436.GSR = "ENABLED";
    FD1P3IX data_buffer__i435 (.D(\data_buffer[427] ), .SP(clk_c_enable_659), 
            .CD(n26795), .CK(clk_c), .Q(\data_buffer[435] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i435.GSR = "ENABLED";
    FD1P3IX data_buffer__i434 (.D(\data_buffer[426] ), .SP(clk_c_enable_659), 
            .CD(n26795), .CK(clk_c), .Q(\data_buffer[434] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i434.GSR = "ENABLED";
    FD1P3IX data_buffer__i433 (.D(\data_buffer[425] ), .SP(clk_c_enable_659), 
            .CD(n26795), .CK(clk_c), .Q(\data_buffer[433] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i433.GSR = "ENABLED";
    FD1P3IX data_buffer__i426 (.D(\data_buffer[418] ), .SP(clk_c_enable_659), 
            .CD(n26795), .CK(clk_c), .Q(\data_buffer[426] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i426.GSR = "ENABLED";
    FD1P3IX data_buffer__i425 (.D(\data_buffer[417] ), .SP(clk_c_enable_659), 
            .CD(n26795), .CK(clk_c), .Q(\data_buffer[425] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i425.GSR = "ENABLED";
    FD1P3IX data_buffer__i424 (.D(\data_buffer[416] ), .SP(clk_c_enable_659), 
            .CD(n26795), .CK(clk_c), .Q(\data_buffer[424] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i424.GSR = "ENABLED";
    FD1P3IX data_buffer__i420 (.D(\data_buffer[412] ), .SP(clk_c_enable_659), 
            .CD(n26795), .CK(clk_c), .Q(\data_buffer[420] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i420.GSR = "ENABLED";
    FD1P3IX data_buffer__i419 (.D(\data_buffer[411] ), .SP(clk_c_enable_659), 
            .CD(n26795), .CK(clk_c), .Q(\data_buffer[419] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i419.GSR = "ENABLED";
    FD1P3IX data_buffer__i418 (.D(\data_buffer[410] ), .SP(clk_c_enable_659), 
            .CD(n26795), .CK(clk_c), .Q(\data_buffer[418] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i418.GSR = "ENABLED";
    FD1P3IX data_buffer__i417 (.D(\data_buffer[409] ), .SP(clk_c_enable_659), 
            .CD(n26795), .CK(clk_c), .Q(\data_buffer[417] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i417.GSR = "ENABLED";
    FD1P3IX data_buffer__i416 (.D(\data_buffer[408] ), .SP(clk_c_enable_659), 
            .CD(n26795), .CK(clk_c), .Q(\data_buffer[416] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i416.GSR = "ENABLED";
    FD1P3IX data_buffer__i412 (.D(\data_buffer[404] ), .SP(clk_c_enable_659), 
            .CD(n26795), .CK(clk_c), .Q(\data_buffer[412] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i412.GSR = "ENABLED";
    FD1P3IX data_buffer__i411 (.D(\data_buffer[403] ), .SP(clk_c_enable_659), 
            .CD(n26795), .CK(clk_c), .Q(\data_buffer[411] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i411.GSR = "ENABLED";
    FD1P3IX data_buffer__i410 (.D(\data_buffer[402] ), .SP(clk_c_enable_659), 
            .CD(n26795), .CK(clk_c), .Q(\data_buffer[410] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i410.GSR = "ENABLED";
    FD1P3IX data_buffer__i409 (.D(\data_buffer[401] ), .SP(clk_c_enable_659), 
            .CD(n26795), .CK(clk_c), .Q(\data_buffer[409] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i409.GSR = "ENABLED";
    FD1P3IX data_buffer__i408 (.D(\data_buffer[400] ), .SP(clk_c_enable_659), 
            .CD(n26795), .CK(clk_c), .Q(\data_buffer[408] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i408.GSR = "ENABLED";
    FD1P3IX data_buffer__i404 (.D(\data_buffer[396] ), .SP(clk_c_enable_659), 
            .CD(n26795), .CK(clk_c), .Q(\data_buffer[404] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i404.GSR = "ENABLED";
    FD1P3IX data_buffer__i403 (.D(\data_buffer[395] ), .SP(clk_c_enable_659), 
            .CD(n26796), .CK(clk_c), .Q(\data_buffer[403] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i403.GSR = "ENABLED";
    FD1P3IX data_buffer__i402 (.D(\data_buffer[394] ), .SP(clk_c_enable_659), 
            .CD(n26796), .CK(clk_c), .Q(\data_buffer[402] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i402.GSR = "ENABLED";
    FD1P3IX data_buffer__i401 (.D(\data_buffer[393] ), .SP(clk_c_enable_659), 
            .CD(n26802), .CK(clk_c), .Q(\data_buffer[401] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i401.GSR = "ENABLED";
    FD1P3IX data_buffer__i400 (.D(\data_buffer[392] ), .SP(clk_c_enable_659), 
            .CD(n26805), .CK(clk_c), .Q(\data_buffer[400] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i400.GSR = "ENABLED";
    FD1P3IX data_buffer__i396 (.D(\data_buffer[388] ), .SP(clk_c_enable_659), 
            .CD(n26796), .CK(clk_c), .Q(\data_buffer[396] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i396.GSR = "ENABLED";
    FD1P3IX data_buffer__i395 (.D(\data_buffer[387] ), .SP(clk_c_enable_659), 
            .CD(n26796), .CK(clk_c), .Q(\data_buffer[395] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i395.GSR = "ENABLED";
    FD1P3IX data_buffer__i394 (.D(\data_buffer[386] ), .SP(clk_c_enable_659), 
            .CD(n26805), .CK(clk_c), .Q(\data_buffer[394] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i394.GSR = "ENABLED";
    FD1P3IX data_buffer__i393 (.D(\data_buffer[385] ), .SP(clk_c_enable_659), 
            .CD(n26796), .CK(clk_c), .Q(\data_buffer[393] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i393.GSR = "ENABLED";
    FD1P3IX data_buffer__i392 (.D(\data_buffer[384] ), .SP(clk_c_enable_659), 
            .CD(n26796), .CK(clk_c), .Q(\data_buffer[392] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i392.GSR = "ENABLED";
    FD1P3IX data_buffer__i388 (.D(\data_buffer[380] ), .SP(clk_c_enable_659), 
            .CD(n26796), .CK(clk_c), .Q(\data_buffer[388] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i388.GSR = "ENABLED";
    FD1P3IX data_buffer__i387 (.D(\data_buffer[379] ), .SP(clk_c_enable_659), 
            .CD(n26796), .CK(clk_c), .Q(\data_buffer[387] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i387.GSR = "ENABLED";
    FD1P3IX data_buffer__i386 (.D(\data_buffer[378] ), .SP(clk_c_enable_659), 
            .CD(n26796), .CK(clk_c), .Q(\data_buffer[386] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i386.GSR = "ENABLED";
    FD1P3IX data_buffer__i385 (.D(\data_buffer[377] ), .SP(clk_c_enable_659), 
            .CD(n26796), .CK(clk_c), .Q(\data_buffer[385] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i385.GSR = "ENABLED";
    FD1P3IX data_buffer__i384 (.D(\data_buffer[376] ), .SP(clk_c_enable_659), 
            .CD(n26796), .CK(clk_c), .Q(\data_buffer[384] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i384.GSR = "ENABLED";
    FD1P3IX data_buffer__i380 (.D(\data_buffer[372] ), .SP(clk_c_enable_659), 
            .CD(n26796), .CK(clk_c), .Q(\data_buffer[380] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i380.GSR = "ENABLED";
    FD1P3IX data_buffer__i379 (.D(\data_buffer[371] ), .SP(clk_c_enable_659), 
            .CD(n26796), .CK(clk_c), .Q(\data_buffer[379] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i379.GSR = "ENABLED";
    FD1P3IX data_buffer__i378 (.D(\data_buffer[370] ), .SP(clk_c_enable_659), 
            .CD(n26796), .CK(clk_c), .Q(\data_buffer[378] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i378.GSR = "ENABLED";
    FD1P3IX data_buffer__i377 (.D(\data_buffer[369] ), .SP(clk_c_enable_659), 
            .CD(n26803), .CK(clk_c), .Q(\data_buffer[377] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i377.GSR = "ENABLED";
    FD1P3IX data_buffer__i376 (.D(\data_buffer[368] ), .SP(clk_c_enable_659), 
            .CD(n26805), .CK(clk_c), .Q(\data_buffer[376] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i376.GSR = "ENABLED";
    FD1P3IX data_buffer__i372 (.D(\data_buffer[364] ), .SP(clk_c_enable_659), 
            .CD(n26796), .CK(clk_c), .Q(\data_buffer[372] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i372.GSR = "ENABLED";
    FD1P3IX data_buffer__i371 (.D(\data_buffer[363] ), .SP(clk_c_enable_659), 
            .CD(n26796), .CK(clk_c), .Q(\data_buffer[371] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i371.GSR = "ENABLED";
    FD1P3IX data_buffer__i370 (.D(\data_buffer[362] ), .SP(clk_c_enable_659), 
            .CD(n26799), .CK(clk_c), .Q(\data_buffer[370] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i370.GSR = "ENABLED";
    FD1P3IX data_buffer__i369 (.D(\data_buffer[361] ), .SP(clk_c_enable_659), 
            .CD(n26805), .CK(clk_c), .Q(\data_buffer[369] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i369.GSR = "ENABLED";
    FD1P3IX data_buffer__i368 (.D(\data_buffer[360] ), .SP(clk_c_enable_659), 
            .CD(n26803), .CK(clk_c), .Q(\data_buffer[368] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i368.GSR = "ENABLED";
    FD1P3IX data_buffer__i364 (.D(\data_buffer[356] ), .SP(clk_c_enable_659), 
            .CD(n26805), .CK(clk_c), .Q(\data_buffer[364] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i364.GSR = "ENABLED";
    FD1P3IX data_buffer__i363 (.D(\data_buffer[355] ), .SP(clk_c_enable_659), 
            .CD(n26803), .CK(clk_c), .Q(\data_buffer[363] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i363.GSR = "ENABLED";
    FD1P3IX data_buffer__i362 (.D(\data_buffer[354] ), .SP(clk_c_enable_659), 
            .CD(n26805), .CK(clk_c), .Q(\data_buffer[362] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i362.GSR = "ENABLED";
    FD1P3IX data_buffer__i361 (.D(\data_buffer[353] ), .SP(clk_c_enable_659), 
            .CD(n26796), .CK(clk_c), .Q(\data_buffer[361] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i361.GSR = "ENABLED";
    FD1P3IX data_buffer__i360 (.D(\data_buffer[352] ), .SP(clk_c_enable_659), 
            .CD(n26803), .CK(clk_c), .Q(\data_buffer[360] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i360.GSR = "ENABLED";
    FD1P3IX data_buffer__i356 (.D(\data_buffer[348] ), .SP(clk_c_enable_659), 
            .CD(n26805), .CK(clk_c), .Q(\data_buffer[356] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i356.GSR = "ENABLED";
    FD1P3IX data_buffer__i355 (.D(\data_buffer[347] ), .SP(clk_c_enable_659), 
            .CD(n26803), .CK(clk_c), .Q(\data_buffer[355] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i355.GSR = "ENABLED";
    FD1P3IX data_buffer__i354 (.D(\data_buffer[346] ), .SP(clk_c_enable_659), 
            .CD(n26796), .CK(clk_c), .Q(\data_buffer[354] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i354.GSR = "ENABLED";
    FD1P3IX data_buffer__i353 (.D(\data_buffer[345] ), .SP(clk_c_enable_659), 
            .CD(n26796), .CK(clk_c), .Q(\data_buffer[353] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i353.GSR = "ENABLED";
    FD1P3IX data_buffer__i352 (.D(\data_buffer[344] ), .SP(clk_c_enable_659), 
            .CD(n26796), .CK(clk_c), .Q(\data_buffer[352] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i352.GSR = "ENABLED";
    FD1P3IX data_buffer__i348 (.D(\data_buffer[340] ), .SP(clk_c_enable_659), 
            .CD(n26796), .CK(clk_c), .Q(\data_buffer[348] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i348.GSR = "ENABLED";
    FD1P3IX data_buffer__i347 (.D(\data_buffer[339] ), .SP(clk_c_enable_659), 
            .CD(n26796), .CK(clk_c), .Q(\data_buffer[347] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i347.GSR = "ENABLED";
    FD1P3IX data_buffer__i346 (.D(\data_buffer[338] ), .SP(clk_c_enable_659), 
            .CD(n26796), .CK(clk_c), .Q(\data_buffer[346] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i346.GSR = "ENABLED";
    FD1P3IX data_buffer__i345 (.D(\data_buffer[337] ), .SP(clk_c_enable_659), 
            .CD(n26796), .CK(clk_c), .Q(\data_buffer[345] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i345.GSR = "ENABLED";
    FD1P3IX data_buffer__i344 (.D(\data_buffer[336] ), .SP(clk_c_enable_659), 
            .CD(n26796), .CK(clk_c), .Q(\data_buffer[344] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i344.GSR = "ENABLED";
    FD1P3IX data_buffer__i340 (.D(\data_buffer[332] ), .SP(clk_c_enable_659), 
            .CD(n26796), .CK(clk_c), .Q(\data_buffer[340] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i340.GSR = "ENABLED";
    FD1P3IX data_buffer__i339 (.D(\data_buffer[331] ), .SP(clk_c_enable_659), 
            .CD(n26796), .CK(clk_c), .Q(\data_buffer[339] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i339.GSR = "ENABLED";
    FD1P3IX data_buffer__i338 (.D(\data_buffer[330] ), .SP(clk_c_enable_659), 
            .CD(n26796), .CK(clk_c), .Q(\data_buffer[338] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i338.GSR = "ENABLED";
    FD1P3IX data_buffer__i337 (.D(\data_buffer[329] ), .SP(clk_c_enable_659), 
            .CD(n26796), .CK(clk_c), .Q(\data_buffer[337] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i337.GSR = "ENABLED";
    FD1P3IX data_buffer__i336 (.D(\data_buffer[328] ), .SP(clk_c_enable_659), 
            .CD(n26796), .CK(clk_c), .Q(\data_buffer[336] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i336.GSR = "ENABLED";
    FD1P3IX data_buffer__i332 (.D(\data_buffer[324] ), .SP(clk_c_enable_659), 
            .CD(n26796), .CK(clk_c), .Q(\data_buffer[332] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i332.GSR = "ENABLED";
    FD1P3IX data_buffer__i331 (.D(\data_buffer[323] ), .SP(clk_c_enable_659), 
            .CD(n26796), .CK(clk_c), .Q(\data_buffer[331] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i331.GSR = "ENABLED";
    FD1P3IX data_buffer__i330 (.D(\data_buffer[322] ), .SP(clk_c_enable_659), 
            .CD(n26796), .CK(clk_c), .Q(\data_buffer[330] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i330.GSR = "ENABLED";
    FD1P3IX data_buffer__i329 (.D(\data_buffer[321] ), .SP(clk_c_enable_659), 
            .CD(n26796), .CK(clk_c), .Q(\data_buffer[329] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i329.GSR = "ENABLED";
    FD1P3IX data_buffer__i328 (.D(\data_buffer[320] ), .SP(clk_c_enable_659), 
            .CD(n26796), .CK(clk_c), .Q(\data_buffer[328] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i328.GSR = "ENABLED";
    FD1P3IX data_buffer__i324 (.D(\data_buffer[316] ), .SP(clk_c_enable_659), 
            .CD(n26796), .CK(clk_c), .Q(\data_buffer[324] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i324.GSR = "ENABLED";
    FD1P3IX data_buffer__i323 (.D(\data_buffer[315] ), .SP(clk_c_enable_659), 
            .CD(n26796), .CK(clk_c), .Q(\data_buffer[323] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i323.GSR = "ENABLED";
    FD1P3IX data_buffer__i322 (.D(\data_buffer[314] ), .SP(clk_c_enable_659), 
            .CD(n26796), .CK(clk_c), .Q(\data_buffer[322] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i322.GSR = "ENABLED";
    FD1P3IX data_buffer__i321 (.D(\data_buffer[313] ), .SP(clk_c_enable_659), 
            .CD(n26796), .CK(clk_c), .Q(\data_buffer[321] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i321.GSR = "ENABLED";
    FD1P3IX data_buffer__i320 (.D(\data_buffer[312] ), .SP(clk_c_enable_659), 
            .CD(n26796), .CK(clk_c), .Q(\data_buffer[320] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i320.GSR = "ENABLED";
    FD1P3IX data_buffer__i316 (.D(\data_buffer[308] ), .SP(clk_c_enable_659), 
            .CD(n26797), .CK(clk_c), .Q(\data_buffer[316] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i316.GSR = "ENABLED";
    FD1P3IX data_buffer__i315 (.D(\data_buffer[307] ), .SP(clk_c_enable_659), 
            .CD(n26796), .CK(clk_c), .Q(\data_buffer[315] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i315.GSR = "ENABLED";
    FD1P3IX data_buffer__i314 (.D(\data_buffer[306] ), .SP(clk_c_enable_659), 
            .CD(n26796), .CK(clk_c), .Q(\data_buffer[314] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i314.GSR = "ENABLED";
    FD1P3IX data_buffer__i313 (.D(\data_buffer[305] ), .SP(clk_c_enable_659), 
            .CD(n26796), .CK(clk_c), .Q(\data_buffer[313] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i313.GSR = "ENABLED";
    FD1P3IX data_buffer__i312 (.D(\data_buffer[304] ), .SP(clk_c_enable_659), 
            .CD(n26796), .CK(clk_c), .Q(\data_buffer[312] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i312.GSR = "ENABLED";
    FD1P3IX data_buffer__i308 (.D(\data_buffer[300] ), .SP(clk_c_enable_659), 
            .CD(n26796), .CK(clk_c), .Q(\data_buffer[308] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i308.GSR = "ENABLED";
    FD1P3IX data_buffer__i307 (.D(\data_buffer[299] ), .SP(clk_c_enable_659), 
            .CD(n26796), .CK(clk_c), .Q(\data_buffer[307] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i307.GSR = "ENABLED";
    FD1P3IX data_buffer__i306 (.D(\data_buffer[298] ), .SP(clk_c_enable_659), 
            .CD(n26805), .CK(clk_c), .Q(\data_buffer[306] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i306.GSR = "ENABLED";
    FD1P3IX data_buffer__i305 (.D(\data_buffer[297] ), .SP(clk_c_enable_659), 
            .CD(n26796), .CK(clk_c), .Q(\data_buffer[305] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i305.GSR = "ENABLED";
    FD1P3IX data_buffer__i304 (.D(\data_buffer[296] ), .SP(clk_c_enable_659), 
            .CD(n26805), .CK(clk_c), .Q(\data_buffer[304] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i304.GSR = "ENABLED";
    FD1P3IX data_buffer__i300 (.D(\data_buffer[292] ), .SP(clk_c_enable_659), 
            .CD(n26799), .CK(clk_c), .Q(\data_buffer[300] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i300.GSR = "ENABLED";
    FD1P3IX data_buffer__i299 (.D(\data_buffer[291] ), .SP(clk_c_enable_659), 
            .CD(n26797), .CK(clk_c), .Q(\data_buffer[299] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i299.GSR = "ENABLED";
    FD1P3IX data_buffer__i298 (.D(\data_buffer[290] ), .SP(clk_c_enable_659), 
            .CD(n26797), .CK(clk_c), .Q(\data_buffer[298] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i298.GSR = "ENABLED";
    FD1P3IX data_buffer__i297 (.D(\data_buffer[289] ), .SP(clk_c_enable_659), 
            .CD(n26799), .CK(clk_c), .Q(\data_buffer[297] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i297.GSR = "ENABLED";
    FD1P3IX data_buffer__i296 (.D(\data_buffer[288] ), .SP(clk_c_enable_659), 
            .CD(n26797), .CK(clk_c), .Q(\data_buffer[296] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i296.GSR = "ENABLED";
    FD1P3IX data_buffer__i292 (.D(\data_buffer[284] ), .SP(clk_c_enable_659), 
            .CD(n26803), .CK(clk_c), .Q(\data_buffer[292] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i292.GSR = "ENABLED";
    FD1P3IX data_buffer__i291 (.D(\data_buffer[283] ), .SP(clk_c_enable_659), 
            .CD(n26799), .CK(clk_c), .Q(\data_buffer[291] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i291.GSR = "ENABLED";
    FD1P3IX data_buffer__i290 (.D(\data_buffer[282] ), .SP(clk_c_enable_659), 
            .CD(n26805), .CK(clk_c), .Q(\data_buffer[290] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i290.GSR = "ENABLED";
    FD1P3IX data_buffer__i289 (.D(\data_buffer[281] ), .SP(clk_c_enable_659), 
            .CD(n26799), .CK(clk_c), .Q(\data_buffer[289] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i289.GSR = "ENABLED";
    FD1P3IX data_buffer__i288 (.D(\data_buffer[280] ), .SP(clk_c_enable_659), 
            .CD(n26800), .CK(clk_c), .Q(\data_buffer[288] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i288.GSR = "ENABLED";
    FD1P3IX data_buffer__i284 (.D(\data_buffer[276] ), .SP(clk_c_enable_659), 
            .CD(n26803), .CK(clk_c), .Q(\data_buffer[284] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i284.GSR = "ENABLED";
    FD1P3IX data_buffer__i283 (.D(\data_buffer[275] ), .SP(clk_c_enable_659), 
            .CD(n26799), .CK(clk_c), .Q(\data_buffer[283] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i283.GSR = "ENABLED";
    FD1P3IX data_buffer__i282 (.D(\data_buffer[274] ), .SP(clk_c_enable_659), 
            .CD(n26802), .CK(clk_c), .Q(\data_buffer[282] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i282.GSR = "ENABLED";
    FD1P3IX data_buffer__i281 (.D(\data_buffer[273] ), .SP(clk_c_enable_659), 
            .CD(n26803), .CK(clk_c), .Q(\data_buffer[281] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i281.GSR = "ENABLED";
    FD1P3IX data_buffer__i280 (.D(\data_buffer[272] ), .SP(clk_c_enable_659), 
            .CD(n26802), .CK(clk_c), .Q(\data_buffer[280] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i280.GSR = "ENABLED";
    FD1P3IX data_buffer__i276 (.D(\data_buffer[268] ), .SP(clk_c_enable_659), 
            .CD(n26805), .CK(clk_c), .Q(\data_buffer[276] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i276.GSR = "ENABLED";
    FD1P3IX data_buffer__i275 (.D(\data_buffer[267] ), .SP(clk_c_enable_659), 
            .CD(n26797), .CK(clk_c), .Q(\data_buffer[275] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i275.GSR = "ENABLED";
    FD1P3IX data_buffer__i274 (.D(\data_buffer[266] ), .SP(clk_c_enable_659), 
            .CD(n26797), .CK(clk_c), .Q(\data_buffer[274] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i274.GSR = "ENABLED";
    FD1P3IX data_buffer__i273 (.D(\data_buffer[265] ), .SP(clk_c_enable_659), 
            .CD(n26805), .CK(clk_c), .Q(\data_buffer[273] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i273.GSR = "ENABLED";
    FD1P3IX data_buffer__i272 (.D(\data_buffer[264] ), .SP(clk_c_enable_659), 
            .CD(n26805), .CK(clk_c), .Q(\data_buffer[272] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i272.GSR = "ENABLED";
    FD1P3IX data_buffer__i268 (.D(\data_buffer[260] ), .SP(clk_c_enable_659), 
            .CD(n26803), .CK(clk_c), .Q(\data_buffer[268] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i268.GSR = "ENABLED";
    FD1P3IX data_buffer__i267 (.D(\data_buffer[259] ), .SP(clk_c_enable_659), 
            .CD(n26805), .CK(clk_c), .Q(\data_buffer[267] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i267.GSR = "ENABLED";
    FD1P3IX data_buffer__i266 (.D(\data_buffer[258] ), .SP(clk_c_enable_659), 
            .CD(n26799), .CK(clk_c), .Q(\data_buffer[266] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i266.GSR = "ENABLED";
    FD1P3IX data_buffer__i265 (.D(\data_buffer[257] ), .SP(clk_c_enable_659), 
            .CD(n26797), .CK(clk_c), .Q(\data_buffer[265] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i265.GSR = "ENABLED";
    FD1P3IX data_buffer__i264 (.D(\data_buffer[256] ), .SP(clk_c_enable_659), 
            .CD(n26805), .CK(clk_c), .Q(\data_buffer[264] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i264.GSR = "ENABLED";
    FD1P3IX data_buffer__i260 (.D(\data_buffer[252] ), .SP(clk_c_enable_659), 
            .CD(n26797), .CK(clk_c), .Q(\data_buffer[260] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i260.GSR = "ENABLED";
    FD1P3IX data_buffer__i259 (.D(\data_buffer[251] ), .SP(clk_c_enable_659), 
            .CD(n26797), .CK(clk_c), .Q(\data_buffer[259] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i259.GSR = "ENABLED";
    FD1P3IX data_buffer__i258 (.D(\data_buffer[250] ), .SP(clk_c_enable_659), 
            .CD(n26803), .CK(clk_c), .Q(\data_buffer[258] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i258.GSR = "ENABLED";
    FD1P3IX data_buffer__i257 (.D(\data_buffer[249] ), .SP(clk_c_enable_659), 
            .CD(n26805), .CK(clk_c), .Q(\data_buffer[257] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i257.GSR = "ENABLED";
    FD1P3IX data_buffer__i256 (.D(\data_buffer[248] ), .SP(clk_c_enable_659), 
            .CD(n26799), .CK(clk_c), .Q(\data_buffer[256] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i256.GSR = "ENABLED";
    FD1P3IX data_buffer__i252 (.D(\data_buffer[244] ), .SP(clk_c_enable_659), 
            .CD(n26797), .CK(clk_c), .Q(\data_buffer[252] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i252.GSR = "ENABLED";
    FD1P3IX data_buffer__i251 (.D(\data_buffer[243] ), .SP(clk_c_enable_659), 
            .CD(n26800), .CK(clk_c), .Q(\data_buffer[251] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i251.GSR = "ENABLED";
    FD1P3IX data_buffer__i250 (.D(\data_buffer[242] ), .SP(clk_c_enable_659), 
            .CD(n26800), .CK(clk_c), .Q(\data_buffer[250] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i250.GSR = "ENABLED";
    FD1P3IX data_buffer__i249 (.D(\data_buffer[241] ), .SP(clk_c_enable_659), 
            .CD(n26800), .CK(clk_c), .Q(\data_buffer[249] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i249.GSR = "ENABLED";
    FD1P3IX data_buffer__i248 (.D(\data_buffer[240] ), .SP(clk_c_enable_659), 
            .CD(n26797), .CK(clk_c), .Q(\data_buffer[248] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i248.GSR = "ENABLED";
    FD1P3IX data_buffer__i244 (.D(\data_buffer[236] ), .SP(clk_c_enable_659), 
            .CD(n26800), .CK(clk_c), .Q(\data_buffer[244] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i244.GSR = "ENABLED";
    FD1P3IX data_buffer__i243 (.D(\data_buffer[235] ), .SP(clk_c_enable_659), 
            .CD(n26797), .CK(clk_c), .Q(\data_buffer[243] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i243.GSR = "ENABLED";
    FD1P3IX data_buffer__i242 (.D(\data_buffer[234] ), .SP(clk_c_enable_659), 
            .CD(n26800), .CK(clk_c), .Q(\data_buffer[242] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i242.GSR = "ENABLED";
    FD1P3IX data_buffer__i241 (.D(\data_buffer[233] ), .SP(clk_c_enable_659), 
            .CD(n26800), .CK(clk_c), .Q(\data_buffer[241] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i241.GSR = "ENABLED";
    FD1P3IX data_buffer__i240 (.D(\data_buffer[232] ), .SP(clk_c_enable_659), 
            .CD(n26797), .CK(clk_c), .Q(\data_buffer[240] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i240.GSR = "ENABLED";
    FD1P3IX data_buffer__i236 (.D(\data_buffer[228] ), .SP(clk_c_enable_659), 
            .CD(n26797), .CK(clk_c), .Q(\data_buffer[236] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i236.GSR = "ENABLED";
    FD1P3IX data_buffer__i235 (.D(\data_buffer[227] ), .SP(clk_c_enable_659), 
            .CD(n26797), .CK(clk_c), .Q(\data_buffer[235] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i235.GSR = "ENABLED";
    FD1P3IX data_buffer__i234 (.D(\data_buffer[226] ), .SP(clk_c_enable_659), 
            .CD(n26800), .CK(clk_c), .Q(\data_buffer[234] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i234.GSR = "ENABLED";
    FD1P3IX data_buffer__i233 (.D(\data_buffer[225] ), .SP(clk_c_enable_659), 
            .CD(n26797), .CK(clk_c), .Q(\data_buffer[233] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i233.GSR = "ENABLED";
    FD1P3IX data_buffer__i232 (.D(\data_buffer[224] ), .SP(clk_c_enable_659), 
            .CD(n26797), .CK(clk_c), .Q(\data_buffer[232] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i232.GSR = "ENABLED";
    FD1P3IX data_buffer__i228 (.D(\data_buffer[220] ), .SP(clk_c_enable_659), 
            .CD(n26800), .CK(clk_c), .Q(\data_buffer[228] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i228.GSR = "ENABLED";
    FD1P3IX data_buffer__i227 (.D(\data_buffer[219] ), .SP(clk_c_enable_659), 
            .CD(n26800), .CK(clk_c), .Q(\data_buffer[227] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i227.GSR = "ENABLED";
    FD1P3IX data_buffer__i226 (.D(\data_buffer[218] ), .SP(clk_c_enable_659), 
            .CD(n26800), .CK(clk_c), .Q(\data_buffer[226] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i226.GSR = "ENABLED";
    FD1P3IX data_buffer__i225 (.D(\data_buffer[217] ), .SP(clk_c_enable_659), 
            .CD(n26797), .CK(clk_c), .Q(\data_buffer[225] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i225.GSR = "ENABLED";
    FD1P3IX rx_done_64_rep_496 (.D(n26780), .SP(rx_done_N_2858), .CD(n26794), 
            .CK(clk_c), .Q(n26793)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(101[10] 104[25])
    defparam rx_done_64_rep_496.GSR = "ENABLED";
    FD1P3IX data_buffer__i224 (.D(\data_buffer[216] ), .SP(clk_c_enable_659), 
            .CD(n26800), .CK(clk_c), .Q(\data_buffer[224] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i224.GSR = "ENABLED";
    FD1P3IX data_buffer__i220 (.D(\data_buffer[212] ), .SP(clk_c_enable_659), 
            .CD(n26800), .CK(clk_c), .Q(\data_buffer[220] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i220.GSR = "ENABLED";
    FD1P3IX data_buffer__i219 (.D(\data_buffer[211] ), .SP(clk_c_enable_659), 
            .CD(n26800), .CK(clk_c), .Q(\data_buffer[219] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i219.GSR = "ENABLED";
    FD1P3IX data_buffer__i218 (.D(\data_buffer[210] ), .SP(clk_c_enable_659), 
            .CD(n26797), .CK(clk_c), .Q(\data_buffer[218] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i218.GSR = "ENABLED";
    FD1P3IX data_buffer__i217 (.D(\data_buffer[209] ), .SP(clk_c_enable_659), 
            .CD(n26800), .CK(clk_c), .Q(\data_buffer[217] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i217.GSR = "ENABLED";
    FD1P3IX data_buffer__i216 (.D(\data_buffer[208] ), .SP(clk_c_enable_659), 
            .CD(n26800), .CK(clk_c), .Q(\data_buffer[216] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i216.GSR = "ENABLED";
    FD1P3IX data_buffer__i212 (.D(\data_buffer[204] ), .SP(clk_c_enable_659), 
            .CD(n26797), .CK(clk_c), .Q(\data_buffer[212] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i212.GSR = "ENABLED";
    FD1P3IX data_buffer__i211 (.D(\data_buffer[203] ), .SP(clk_c_enable_659), 
            .CD(n26800), .CK(clk_c), .Q(\data_buffer[211] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i211.GSR = "ENABLED";
    FD1P3IX data_buffer__i210 (.D(\data_buffer[202] ), .SP(clk_c_enable_659), 
            .CD(n26800), .CK(clk_c), .Q(\data_buffer[210] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i210.GSR = "ENABLED";
    FD1P3IX data_buffer__i209 (.D(\data_buffer[201] ), .SP(clk_c_enable_659), 
            .CD(n26800), .CK(clk_c), .Q(\data_buffer[209] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i209.GSR = "ENABLED";
    FD1P3IX data_buffer__i208 (.D(\data_buffer[200] ), .SP(clk_c_enable_659), 
            .CD(n26800), .CK(clk_c), .Q(\data_buffer[208] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i208.GSR = "ENABLED";
    FD1P3IX data_buffer__i204 (.D(\data_buffer[196] ), .SP(clk_c_enable_659), 
            .CD(n26797), .CK(clk_c), .Q(\data_buffer[204] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i204.GSR = "ENABLED";
    FD1P3IX data_buffer__i203 (.D(\data_buffer[195] ), .SP(clk_c_enable_659), 
            .CD(n26803), .CK(clk_c), .Q(\data_buffer[203] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i203.GSR = "ENABLED";
    FD1P3IX data_buffer__i202 (.D(\data_buffer[194] ), .SP(clk_c_enable_659), 
            .CD(n26800), .CK(clk_c), .Q(\data_buffer[202] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i202.GSR = "ENABLED";
    FD1P3IX data_buffer__i201 (.D(\data_buffer[193] ), .SP(clk_c_enable_659), 
            .CD(n26805), .CK(clk_c), .Q(\data_buffer[201] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i201.GSR = "ENABLED";
    FD1P3IX data_buffer__i200 (.D(\data_buffer[192] ), .SP(clk_c_enable_659), 
            .CD(n26800), .CK(clk_c), .Q(\data_buffer[200] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i200.GSR = "ENABLED";
    FD1P3IX data_buffer__i196 (.D(\data_buffer[188] ), .SP(clk_c_enable_659), 
            .CD(n26800), .CK(clk_c), .Q(\data_buffer[196] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i196.GSR = "ENABLED";
    FD1P3IX data_buffer__i195 (.D(\data_buffer[187] ), .SP(clk_c_enable_659), 
            .CD(n26802), .CK(clk_c), .Q(\data_buffer[195] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i195.GSR = "ENABLED";
    FD1P3IX data_buffer__i178 (.D(\data_buffer[170] ), .SP(clk_c_enable_659), 
            .CD(n26800), .CK(clk_c), .Q(\data_buffer[178] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i178.GSR = "ENABLED";
    FD1P3IX data_buffer__i179 (.D(\data_buffer[171] ), .SP(clk_c_enable_659), 
            .CD(n26800), .CK(clk_c), .Q(\data_buffer[179] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i179.GSR = "ENABLED";
    FD1P3IX data_buffer__i180 (.D(\data_buffer[172] ), .SP(clk_c_enable_659), 
            .CD(n26800), .CK(clk_c), .Q(\data_buffer[180] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i180.GSR = "ENABLED";
    FD1P3IX data_buffer__i184 (.D(\data_buffer[176] ), .SP(clk_c_enable_659), 
            .CD(n26800), .CK(clk_c), .Q(\data_buffer[184] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i184.GSR = "ENABLED";
    FD1P3IX data_buffer__i185 (.D(\data_buffer[177] ), .SP(clk_c_enable_659), 
            .CD(n26800), .CK(clk_c), .Q(\data_buffer[185] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i185.GSR = "ENABLED";
    FD1P3IX data_buffer__i186 (.D(\data_buffer[178] ), .SP(clk_c_enable_659), 
            .CD(n26803), .CK(clk_c), .Q(\data_buffer[186] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i186.GSR = "ENABLED";
    FD1P3IX data_buffer__i187 (.D(\data_buffer[179] ), .SP(clk_c_enable_659), 
            .CD(n26800), .CK(clk_c), .Q(\data_buffer[187] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i187.GSR = "ENABLED";
    FD1P3IX data_buffer__i188 (.D(\data_buffer[180] ), .SP(clk_c_enable_659), 
            .CD(n26805), .CK(clk_c), .Q(\data_buffer[188] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i188.GSR = "ENABLED";
    FD1P3IX data_buffer__i192 (.D(\data_buffer[184] ), .SP(clk_c_enable_659), 
            .CD(n26800), .CK(clk_c), .Q(\data_buffer[192] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i192.GSR = "ENABLED";
    FD1P3IX data_buffer__i193 (.D(\data_buffer[185] ), .SP(clk_c_enable_659), 
            .CD(n26800), .CK(clk_c), .Q(\data_buffer[193] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i193.GSR = "ENABLED";
    FD1P3IX data_buffer__i194 (.D(\data_buffer[186] ), .SP(clk_c_enable_659), 
            .CD(n26800), .CK(clk_c), .Q(\data_buffer[194] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i194.GSR = "ENABLED";
    FD1P3IX data_buffer__i177 (.D(\data_buffer[169] ), .SP(clk_c_enable_659), 
            .CD(n26800), .CK(clk_c), .Q(\data_buffer[177] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i177.GSR = "ENABLED";
    FD1P3IX data_buffer__i176 (.D(\data_buffer[168] ), .SP(clk_c_enable_659), 
            .CD(n26800), .CK(clk_c), .Q(\data_buffer[176] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i176.GSR = "ENABLED";
    FD1P3IX data_buffer__i172 (.D(\data_buffer[164] ), .SP(clk_c_enable_659), 
            .CD(n26803), .CK(clk_c), .Q(\data_buffer[172] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i172.GSR = "ENABLED";
    FD1P3IX data_buffer__i171 (.D(\data_buffer[163] ), .SP(clk_c_enable_659), 
            .CD(n26800), .CK(clk_c), .Q(\data_buffer[171] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i171.GSR = "ENABLED";
    FD1P3IX data_buffer__i170 (.D(\data_buffer[162] ), .SP(clk_c_enable_659), 
            .CD(n26805), .CK(clk_c), .Q(\data_buffer[170] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i170.GSR = "ENABLED";
    FD1P3IX data_buffer__i169 (.D(\data_buffer[161] ), .SP(clk_c_enable_659), 
            .CD(n26797), .CK(clk_c), .Q(\data_buffer[169] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i169.GSR = "ENABLED";
    FD1P3IX data_buffer__i168 (.D(\data_buffer[160] ), .SP(clk_c_enable_659), 
            .CD(n26800), .CK(clk_c), .Q(\data_buffer[168] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i168.GSR = "ENABLED";
    FD1P3IX data_buffer__i164 (.D(\data_buffer[156] ), .SP(clk_c_enable_659), 
            .CD(n26800), .CK(clk_c), .Q(\data_buffer[164] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i164.GSR = "ENABLED";
    FD1P3IX data_buffer__i163 (.D(\data_buffer[155] ), .SP(clk_c_enable_659), 
            .CD(n26800), .CK(clk_c), .Q(\data_buffer[163] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i163.GSR = "ENABLED";
    FD1P3IX data_buffer__i162 (.D(\data_buffer[154] ), .SP(clk_c_enable_659), 
            .CD(n26805), .CK(clk_c), .Q(\data_buffer[162] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i162.GSR = "ENABLED";
    FD1P3IX data_buffer__i161 (.D(\data_buffer[153] ), .SP(clk_c_enable_659), 
            .CD(n26800), .CK(clk_c), .Q(\data_buffer[161] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i161.GSR = "ENABLED";
    FD1P3IX data_buffer__i160 (.D(\data_buffer[152] ), .SP(clk_c_enable_659), 
            .CD(n26800), .CK(clk_c), .Q(\data_buffer[160] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i160.GSR = "ENABLED";
    FD1P3IX data_buffer__i156 (.D(\data_buffer[148] ), .SP(clk_c_enable_659), 
            .CD(n26805), .CK(clk_c), .Q(\data_buffer[156] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i156.GSR = "ENABLED";
    FD1P3IX data_buffer__i155 (.D(\data_buffer[147] ), .SP(clk_c_enable_659), 
            .CD(n26800), .CK(clk_c), .Q(\data_buffer[155] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i155.GSR = "ENABLED";
    FD1P3IX data_buffer__i154 (.D(\data_buffer[146] ), .SP(clk_c_enable_659), 
            .CD(n26800), .CK(clk_c), .Q(\data_buffer[154] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i154.GSR = "ENABLED";
    FD1P3IX data_buffer__i153 (.D(\data_buffer[145] ), .SP(clk_c_enable_659), 
            .CD(n26805), .CK(clk_c), .Q(\data_buffer[153] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i153.GSR = "ENABLED";
    FD1P3IX data_buffer__i152 (.D(\data_buffer[144] ), .SP(clk_c_enable_659), 
            .CD(n26800), .CK(clk_c), .Q(\data_buffer[152] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i152.GSR = "ENABLED";
    FD1P3IX data_buffer__i148 (.D(\data_buffer[140] ), .SP(clk_c_enable_659), 
            .CD(n26800), .CK(clk_c), .Q(\data_buffer[148] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i148.GSR = "ENABLED";
    FD1P3IX data_buffer__i147 (.D(\data_buffer[139] ), .SP(clk_c_enable_659), 
            .CD(n26794), .CK(clk_c), .Q(\data_buffer[147] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i147.GSR = "ENABLED";
    FD1P3IX data_buffer__i146 (.D(\data_buffer[138] ), .SP(clk_c_enable_659), 
            .CD(n26801), .CK(clk_c), .Q(\data_buffer[146] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i146.GSR = "ENABLED";
    FD1P3IX data_buffer__i145 (.D(\data_buffer[137] ), .SP(clk_c_enable_659), 
            .CD(n26797), .CK(clk_c), .Q(\data_buffer[145] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i145.GSR = "ENABLED";
    FD1P3IX data_buffer__i144 (.D(\data_buffer[136] ), .SP(clk_c_enable_659), 
            .CD(n26801), .CK(clk_c), .Q(\data_buffer[144] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i144.GSR = "ENABLED";
    FD1P3IX data_buffer__i140 (.D(\data_buffer[132] ), .SP(clk_c_enable_659), 
            .CD(n26801), .CK(clk_c), .Q(\data_buffer[140] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i140.GSR = "ENABLED";
    FD1P3IX data_buffer__i139 (.D(\data_buffer[131] ), .SP(clk_c_enable_659), 
            .CD(n26801), .CK(clk_c), .Q(\data_buffer[139] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i139.GSR = "ENABLED";
    FD1P3IX data_buffer__i138 (.D(\data_buffer[130] ), .SP(clk_c_enable_659), 
            .CD(n26798), .CK(clk_c), .Q(\data_buffer[138] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i138.GSR = "ENABLED";
    FD1P3IX data_buffer__i137 (.D(\data_buffer[129] ), .SP(clk_c_enable_659), 
            .CD(n26801), .CK(clk_c), .Q(\data_buffer[137] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i137.GSR = "ENABLED";
    FD1P3IX data_buffer__i136 (.D(\data_buffer[128] ), .SP(clk_c_enable_659), 
            .CD(n26802), .CK(clk_c), .Q(\data_buffer[136] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i136.GSR = "ENABLED";
    FD1P3IX data_buffer__i132 (.D(\data_buffer[124] ), .SP(clk_c_enable_659), 
            .CD(n26797), .CK(clk_c), .Q(\data_buffer[132] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i132.GSR = "ENABLED";
    FD1P3IX data_buffer__i131 (.D(\data_buffer[123] ), .SP(clk_c_enable_659), 
            .CD(n26801), .CK(clk_c), .Q(\data_buffer[131] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i131.GSR = "ENABLED";
    FD1P3IX data_buffer__i130 (.D(\data_buffer[122] ), .SP(clk_c_enable_659), 
            .CD(n26802), .CK(clk_c), .Q(\data_buffer[130] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i130.GSR = "ENABLED";
    FD1P3IX data_buffer__i129 (.D(\data_buffer[121] ), .SP(clk_c_enable_659), 
            .CD(n26801), .CK(clk_c), .Q(\data_buffer[129] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i129.GSR = "ENABLED";
    FD1P3IX data_buffer__i128 (.D(\data_buffer[120] ), .SP(clk_c_enable_659), 
            .CD(n26797), .CK(clk_c), .Q(\data_buffer[128] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i128.GSR = "ENABLED";
    FD1P3IX data_buffer__i124 (.D(\data_buffer[116] ), .SP(clk_c_enable_659), 
            .CD(n26797), .CK(clk_c), .Q(\data_buffer[124] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i124.GSR = "ENABLED";
    FD1P3IX data_buffer__i123 (.D(\data_buffer[115] ), .SP(clk_c_enable_659), 
            .CD(n26797), .CK(clk_c), .Q(\data_buffer[123] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i123.GSR = "ENABLED";
    FD1P3IX data_buffer__i122 (.D(\data_buffer[114] ), .SP(clk_c_enable_659), 
            .CD(n26797), .CK(clk_c), .Q(\data_buffer[122] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i122.GSR = "ENABLED";
    FD1P3IX data_buffer__i121 (.D(\data_buffer[113] ), .SP(clk_c_enable_659), 
            .CD(n26801), .CK(clk_c), .Q(\data_buffer[121] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i121.GSR = "ENABLED";
    FD1P3IX data_buffer__i120 (.D(\data_buffer[112] ), .SP(clk_c_enable_659), 
            .CD(n26797), .CK(clk_c), .Q(\data_buffer[120] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i120.GSR = "ENABLED";
    FD1P3IX data_buffer__i116 (.D(\data_buffer[108] ), .SP(clk_c_enable_659), 
            .CD(n26801), .CK(clk_c), .Q(\data_buffer[116] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i116.GSR = "ENABLED";
    FD1P3IX data_buffer__i115 (.D(\data_buffer[107] ), .SP(clk_c_enable_659), 
            .CD(n26798), .CK(clk_c), .Q(\data_buffer[115] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i115.GSR = "ENABLED";
    FD1P3IX data_buffer__i114 (.D(\data_buffer[106] ), .SP(clk_c_enable_659), 
            .CD(n26801), .CK(clk_c), .Q(\data_buffer[114] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i114.GSR = "ENABLED";
    FD1P3IX data_buffer__i113 (.D(\data_buffer[105] ), .SP(clk_c_enable_659), 
            .CD(n26797), .CK(clk_c), .Q(\data_buffer[113] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i113.GSR = "ENABLED";
    FD1P3IX data_buffer__i112 (.D(\data_buffer[104] ), .SP(clk_c_enable_659), 
            .CD(n26801), .CK(clk_c), .Q(\data_buffer[112] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i112.GSR = "ENABLED";
    FD1P3IX data_buffer__i108 (.D(\data_buffer[100] ), .SP(clk_c_enable_659), 
            .CD(n26797), .CK(clk_c), .Q(\data_buffer[108] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i108.GSR = "ENABLED";
    FD1P3IX data_buffer__i107 (.D(\data_buffer[99] ), .SP(clk_c_enable_659), 
            .CD(n26803), .CK(clk_c), .Q(\data_buffer[107] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i107.GSR = "ENABLED";
    FD1P3IX data_buffer__i106 (.D(\data_buffer[98] ), .SP(clk_c_enable_659), 
            .CD(n26805), .CK(clk_c), .Q(\data_buffer[106] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i106.GSR = "ENABLED";
    FD1P3IX data_buffer__i105 (.D(\data_buffer[97] ), .SP(clk_c_enable_659), 
            .CD(n26797), .CK(clk_c), .Q(\data_buffer[105] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i105.GSR = "ENABLED";
    FD1P3IX data_buffer__i104 (.D(\data_buffer[96] ), .SP(clk_c_enable_659), 
            .CD(n26801), .CK(clk_c), .Q(\data_buffer[104] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i104.GSR = "ENABLED";
    FD1P3IX data_buffer__i100 (.D(\data_buffer[92] ), .SP(clk_c_enable_659), 
            .CD(n26805), .CK(clk_c), .Q(\data_buffer[100] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i100.GSR = "ENABLED";
    FD1P3IX data_buffer__i99 (.D(\data_buffer[91] ), .SP(clk_c_enable_659), 
            .CD(n26802), .CK(clk_c), .Q(\data_buffer[99] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i99.GSR = "ENABLED";
    FD1P3IX data_buffer__i98 (.D(\data_buffer[90] ), .SP(clk_c_enable_659), 
            .CD(n26803), .CK(clk_c), .Q(\data_buffer[98] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i98.GSR = "ENABLED";
    FD1P3IX data_buffer__i97 (.D(\data_buffer[89] ), .SP(clk_c_enable_659), 
            .CD(n26801), .CK(clk_c), .Q(\data_buffer[97] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i97.GSR = "ENABLED";
    FD1P3IX data_buffer__i96 (.D(\data_buffer[88] ), .SP(clk_c_enable_659), 
            .CD(n26801), .CK(clk_c), .Q(\data_buffer[96] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i96.GSR = "ENABLED";
    FD1P3IX data_buffer__i92 (.D(\data_buffer[84] ), .SP(clk_c_enable_659), 
            .CD(n26805), .CK(clk_c), .Q(\data_buffer[92] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i92.GSR = "ENABLED";
    FD1P3IX data_buffer__i91 (.D(\data_buffer[83] ), .SP(clk_c_enable_659), 
            .CD(n26797), .CK(clk_c), .Q(\data_buffer[91] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i91.GSR = "ENABLED";
    FD1P3IX data_buffer__i90 (.D(\data_buffer[82] ), .SP(clk_c_enable_659), 
            .CD(n26801), .CK(clk_c), .Q(\data_buffer[90] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i90.GSR = "ENABLED";
    FD1P3IX data_buffer__i89 (.D(\data_buffer[81] ), .SP(clk_c_enable_659), 
            .CD(n26801), .CK(clk_c), .Q(\data_buffer[89] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i89.GSR = "ENABLED";
    FD1P3IX data_buffer__i88 (.D(\data_buffer[80] ), .SP(clk_c_enable_659), 
            .CD(n26802), .CK(clk_c), .Q(\data_buffer[88] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i88.GSR = "ENABLED";
    FD1P3IX data_buffer__i84 (.D(\data_buffer[76] ), .SP(clk_c_enable_659), 
            .CD(n26797), .CK(clk_c), .Q(\data_buffer[84] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i84.GSR = "ENABLED";
    FD1P3IX data_buffer__i83 (.D(\data_buffer[75] ), .SP(clk_c_enable_659), 
            .CD(n26797), .CK(clk_c), .Q(\data_buffer[83] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i83.GSR = "ENABLED";
    FD1P3IX data_buffer__i82 (.D(\data_buffer[74] ), .SP(clk_c_enable_659), 
            .CD(n26797), .CK(clk_c), .Q(\data_buffer[82] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i82.GSR = "ENABLED";
    FD1P3IX data_buffer__i81 (.D(\data_buffer[73] ), .SP(clk_c_enable_659), 
            .CD(n26801), .CK(clk_c), .Q(\data_buffer[81] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i81.GSR = "ENABLED";
    FD1P3IX data_length__i0 (.D(n78[0]), .SP(clk_c_enable_1399), .CD(n26797), 
            .CK(clk_c), .Q(data_length[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(79[10] 84[43])
    defparam data_length__i0.GSR = "ENABLED";
    FD1P3IX data_buffer__i80 (.D(\data_buffer[72] ), .SP(clk_c_enable_659), 
            .CD(rx_done), .CK(clk_c), .Q(\data_buffer[80] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i80.GSR = "ENABLED";
    FD1P3IX data_buffer__i76 (.D(\data_buffer[68] ), .SP(clk_c_enable_659), 
            .CD(n26801), .CK(clk_c), .Q(\data_buffer[76] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i76.GSR = "ENABLED";
    FD1P3IX data_buffer__i75 (.D(\data_buffer[67] ), .SP(clk_c_enable_659), 
            .CD(n26797), .CK(clk_c), .Q(\data_buffer[75] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i75.GSR = "ENABLED";
    FD1P3IX data_buffer__i74 (.D(\data_buffer[66] ), .SP(clk_c_enable_659), 
            .CD(n26797), .CK(clk_c), .Q(\data_buffer[74] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i74.GSR = "ENABLED";
    FD1P3IX data_buffer__i73 (.D(\data_buffer[65] ), .SP(clk_c_enable_659), 
            .CD(n26801), .CK(clk_c), .Q(\data_buffer[73] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i73.GSR = "ENABLED";
    FD1P3IX data_buffer__i72 (.D(\data_buffer[64] ), .SP(clk_c_enable_659), 
            .CD(n26798), .CK(clk_c), .Q(\data_buffer[72] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i72.GSR = "ENABLED";
    FD1P3IX data_buffer__i68 (.D(\data_buffer[60] ), .SP(clk_c_enable_659), 
            .CD(n26801), .CK(clk_c), .Q(\data_buffer[68] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i68.GSR = "ENABLED";
    FD1P3IX data_buffer__i67 (.D(\data_buffer[59] ), .SP(clk_c_enable_659), 
            .CD(n26801), .CK(clk_c), .Q(\data_buffer[67] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i67.GSR = "ENABLED";
    FD1P3IX data_buffer__i66 (.D(\data_buffer[58] ), .SP(clk_c_enable_659), 
            .CD(n26801), .CK(clk_c), .Q(\data_buffer[66] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i66.GSR = "ENABLED";
    FD1P3IX data_buffer__i65 (.D(\data_buffer[57] ), .SP(clk_c_enable_659), 
            .CD(n26798), .CK(clk_c), .Q(\data_buffer[65] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i65.GSR = "ENABLED";
    FD1P3IX data_buffer__i64 (.D(\data_buffer[56] ), .SP(clk_c_enable_659), 
            .CD(n26798), .CK(clk_c), .Q(\data_buffer[64] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i64.GSR = "ENABLED";
    FD1P3IX data_buffer__i60 (.D(\data_buffer[52] ), .SP(clk_c_enable_659), 
            .CD(n26797), .CK(clk_c), .Q(\data_buffer[60] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i60.GSR = "ENABLED";
    FD1P3IX data_buffer__i59 (.D(\data_buffer[51] ), .SP(clk_c_enable_659), 
            .CD(n26798), .CK(clk_c), .Q(\data_buffer[59] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i59.GSR = "ENABLED";
    FD1P3IX data_buffer__i58 (.D(\data_buffer[50] ), .SP(clk_c_enable_659), 
            .CD(n26798), .CK(clk_c), .Q(\data_buffer[58] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i58.GSR = "ENABLED";
    FD1P3IX data_buffer__i57 (.D(\data_buffer[49] ), .SP(clk_c_enable_659), 
            .CD(n26801), .CK(clk_c), .Q(\data_buffer[57] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i57.GSR = "ENABLED";
    FD1P3IX data_buffer__i56 (.D(\data_buffer[48] ), .SP(clk_c_enable_659), 
            .CD(n26802), .CK(clk_c), .Q(\data_buffer[56] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i56.GSR = "ENABLED";
    FD1P3IX data_buffer__i52 (.D(\data_buffer[44] ), .SP(clk_c_enable_659), 
            .CD(n26801), .CK(clk_c), .Q(\data_buffer[52] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i52.GSR = "ENABLED";
    FD1P3IX data_buffer__i51 (.D(\data_buffer[43] ), .SP(clk_c_enable_659), 
            .CD(n26801), .CK(clk_c), .Q(\data_buffer[51] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i51.GSR = "ENABLED";
    FD1P3IX data_buffer__i50 (.D(\data_buffer[42] ), .SP(clk_c_enable_659), 
            .CD(n26801), .CK(clk_c), .Q(\data_buffer[50] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i50.GSR = "ENABLED";
    FD1P3IX data_buffer__i49 (.D(\data_buffer[41] ), .SP(clk_c_enable_659), 
            .CD(n26801), .CK(clk_c), .Q(\data_buffer[49] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i49.GSR = "ENABLED";
    FD1P3IX data_buffer__i48 (.D(\data_buffer[40] ), .SP(clk_c_enable_659), 
            .CD(n26798), .CK(clk_c), .Q(\data_buffer[48] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i48.GSR = "ENABLED";
    FD1P3IX data_buffer__i44 (.D(\data_buffer[36] ), .SP(clk_c_enable_659), 
            .CD(n26797), .CK(clk_c), .Q(\data_buffer[44] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i44.GSR = "ENABLED";
    FD1P3IX data_buffer__i43 (.D(\data_buffer[35] ), .SP(clk_c_enable_659), 
            .CD(n26798), .CK(clk_c), .Q(\data_buffer[43] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i43.GSR = "ENABLED";
    FD1P3IX data_buffer__i42 (.D(\data_buffer[34] ), .SP(clk_c_enable_659), 
            .CD(n26798), .CK(clk_c), .Q(\data_buffer[42] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i42.GSR = "ENABLED";
    FD1P3IX data_buffer__i41 (.D(\data_buffer[33] ), .SP(clk_c_enable_659), 
            .CD(n26796), .CK(clk_c), .Q(\data_buffer[41] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i41.GSR = "ENABLED";
    FD1P3IX data_buffer__i40 (.D(\data_buffer[32] ), .SP(clk_c_enable_659), 
            .CD(n26798), .CK(clk_c), .Q(\data_buffer[40] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i40.GSR = "ENABLED";
    FD1P3IX data_buffer__i36 (.D(\data_buffer[28] ), .SP(clk_c_enable_659), 
            .CD(n26796), .CK(clk_c), .Q(\data_buffer[36] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i36.GSR = "ENABLED";
    FD1P3IX data_buffer__i35 (.D(\data_buffer[27] ), .SP(clk_c_enable_659), 
            .CD(n26795), .CK(clk_c), .Q(\data_buffer[35] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i35.GSR = "ENABLED";
    FD1P3IX data_buffer__i34 (.D(\data_buffer[26] ), .SP(clk_c_enable_659), 
            .CD(n26798), .CK(clk_c), .Q(\data_buffer[34] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i34.GSR = "ENABLED";
    FD1P3IX data_buffer__i33 (.D(\data_buffer[25] ), .SP(clk_c_enable_659), 
            .CD(n26798), .CK(clk_c), .Q(\data_buffer[33] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i33.GSR = "ENABLED";
    FD1P3IX data_buffer__i32 (.D(\data_buffer[24] ), .SP(clk_c_enable_659), 
            .CD(n26798), .CK(clk_c), .Q(\data_buffer[32] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i32.GSR = "ENABLED";
    FD1P3IX data_buffer__i28 (.D(\data_buffer[20] ), .SP(clk_c_enable_659), 
            .CD(n26798), .CK(clk_c), .Q(\data_buffer[28] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i28.GSR = "ENABLED";
    FD1P3IX data_buffer__i27 (.D(\data_buffer[19] ), .SP(clk_c_enable_659), 
            .CD(n26798), .CK(clk_c), .Q(\data_buffer[27] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i27.GSR = "ENABLED";
    FD1P3IX data_buffer__i26 (.D(\data_buffer[18] ), .SP(clk_c_enable_659), 
            .CD(n26798), .CK(clk_c), .Q(\data_buffer[26] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i26.GSR = "ENABLED";
    FD1P3IX data_buffer__i25 (.D(\data_buffer[17] ), .SP(clk_c_enable_659), 
            .CD(n26798), .CK(clk_c), .Q(\data_buffer[25] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i25.GSR = "ENABLED";
    FD1P3IX data_buffer__i24 (.D(\data_buffer[16] ), .SP(clk_c_enable_659), 
            .CD(n26798), .CK(clk_c), .Q(\data_buffer[24] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i24.GSR = "ENABLED";
    FD1P3IX data_buffer__i20 (.D(\data_buffer[12] ), .SP(clk_c_enable_659), 
            .CD(n26801), .CK(clk_c), .Q(\data_buffer[20] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i20.GSR = "ENABLED";
    FD1P3IX data_buffer__i19 (.D(\data_buffer[11] ), .SP(clk_c_enable_659), 
            .CD(n26798), .CK(clk_c), .Q(\data_buffer[19] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i19.GSR = "ENABLED";
    FD1P3IX data_buffer__i18 (.D(\data_buffer[10] ), .SP(clk_c_enable_659), 
            .CD(n26798), .CK(clk_c), .Q(\data_buffer[18] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i18.GSR = "ENABLED";
    FD1P3IX data_buffer__i17 (.D(\data_buffer[9] ), .SP(clk_c_enable_659), 
            .CD(n26798), .CK(clk_c), .Q(\data_buffer[17] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i17.GSR = "ENABLED";
    FD1P3IX data_buffer__i16 (.D(\data_buffer[8] ), .SP(clk_c_enable_659), 
            .CD(n26798), .CK(clk_c), .Q(\data_buffer[16] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i16.GSR = "ENABLED";
    FD1P3IX data_buffer__i12 (.D(\data_buffer[4] ), .SP(clk_c_enable_659), 
            .CD(n26801), .CK(clk_c), .Q(\data_buffer[12] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i12.GSR = "ENABLED";
    FD1P3IX data_buffer__i11 (.D(\data_buffer[3] ), .SP(clk_c_enable_659), 
            .CD(rx_done), .CK(clk_c), .Q(\data_buffer[11] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i11.GSR = "ENABLED";
    FD1P3IX data_buffer__i10 (.D(\data_buffer[2] ), .SP(clk_c_enable_659), 
            .CD(n26797), .CK(clk_c), .Q(\data_buffer[10] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i10.GSR = "ENABLED";
    FD1P3IX data_buffer__i9 (.D(\data_buffer[1] ), .SP(clk_c_enable_659), 
            .CD(n26802), .CK(clk_c), .Q(\data_buffer[9] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i9.GSR = "ENABLED";
    FD1P3IX data_buffer__i8 (.D(\data_buffer[0] ), .SP(clk_c_enable_659), 
            .CD(n26802), .CK(clk_c), .Q(\data_buffer[8] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i8.GSR = "ENABLED";
    FD1P3IX data_buffer__i4 (.D(rx_data[4]), .SP(clk_c_enable_659), .CD(n26802), 
            .CK(clk_c), .Q(\data_buffer[4] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i4.GSR = "ENABLED";
    FD1P3IX data_buffer__i3 (.D(rx_data[3]), .SP(clk_c_enable_659), .CD(n26798), 
            .CK(clk_c), .Q(\data_buffer[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i3.GSR = "ENABLED";
    FD1P3IX data_buffer__i2 (.D(rx_data[2]), .SP(clk_c_enable_659), .CD(rx_done), 
            .CK(clk_c), .Q(\data_buffer[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i2.GSR = "ENABLED";
    FD1P3IX data_buffer__i1 (.D(rx_data[1]), .SP(clk_c_enable_659), .CD(rx_done), 
            .CK(clk_c), .Q(\data_buffer[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(89[10] 96[8])
    defparam data_buffer__i1.GSR = "ENABLED";
    FD1P3IX rx_done_64_rep_508 (.D(n26780), .SP(rx_done_N_2858), .CD(n26805), 
            .CK(clk_c), .Q(n26805)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(101[10] 104[25])
    defparam rx_done_64_rep_508.GSR = "ENABLED";
    FD1P3IX rx_done_64 (.D(n26780), .SP(rx_done_N_2858), .CD(rx_done), 
            .CK(clk_c), .Q(rx_done)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(101[10] 104[25])
    defparam rx_done_64.GSR = "ENABLED";
    FD1P3IX tx_data_length_i1 (.D(n9394), .SP(tx_done), .CD(flag), .CK(clk_c), 
            .Q(tx_data_length[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(46[10] 49[49])
    defparam tx_data_length_i1.GSR = "ENABLED";
    FD1P3AX tx_data_i1 (.D(tx_data_7__N_1868[1]), .SP(clk_c_enable_1418), 
            .CK(clk_c), .Q(tx_data[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(56[10] 59[42])
    defparam tx_data_i1.GSR = "ENABLED";
    FD1P3AX tx_data_i2 (.D(tx_data_7__N_1868[2]), .SP(clk_c_enable_1418), 
            .CK(clk_c), .Q(tx_data[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(56[10] 59[42])
    defparam tx_data_i2.GSR = "ENABLED";
    FD1P3AX tx_data_i3 (.D(tx_data_7__N_1868[3]), .SP(clk_c_enable_1418), 
            .CK(clk_c), .Q(tx_data[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(56[10] 59[42])
    defparam tx_data_i3.GSR = "ENABLED";
    LUT4 i9269_2_lut (.A(tx_done), .B(flag), .Z(n12084)) /* synthesis lut_function=(!((B)+!A)) */ ;   // g:/fpga/mxo2/system/project/uart_top.v(56[10] 59[42])
    defparam i9269_2_lut.init = 16'h2222;
    CCU2D add_35_11 (.A0(data_length[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n20509), .S0(n78[9]));   // g:/fpga/mxo2/system/project/uart_top.v(84[24:42])
    defparam add_35_11.INIT0 = 16'h5aaa;
    defparam add_35_11.INIT1 = 16'h0000;
    defparam add_35_11.INJECT1_0 = "NO";
    defparam add_35_11.INJECT1_1 = "NO";
    FD1P3IX rx_done_64_rep_507 (.D(n26780), .SP(rx_done_N_2858), .CD(n26804), 
            .CK(clk_c), .Q(n26804)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(101[10] 104[25])
    defparam rx_done_64_rep_507.GSR = "ENABLED";
    CCU2D add_35_9 (.A0(data_length[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(data_length[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n20508), .COUT(n20509), .S0(n78[7]), .S1(n78[8]));   // g:/fpga/mxo2/system/project/uart_top.v(84[24:42])
    defparam add_35_9.INIT0 = 16'h5aaa;
    defparam add_35_9.INIT1 = 16'h5aaa;
    defparam add_35_9.INJECT1_0 = "NO";
    defparam add_35_9.INJECT1_1 = "NO";
    CCU2D add_35_7 (.A0(data_length[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(data_length[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n20507), .COUT(n20508), .S0(n78[5]), .S1(n78[6]));   // g:/fpga/mxo2/system/project/uart_top.v(84[24:42])
    defparam add_35_7.INIT0 = 16'h5aaa;
    defparam add_35_7.INIT1 = 16'h5aaa;
    defparam add_35_7.INJECT1_0 = "NO";
    defparam add_35_7.INJECT1_1 = "NO";
    CCU2D add_35_5 (.A0(data_length[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(data_length[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n20506), .COUT(n20507), .S0(n78[3]), .S1(n78[4]));   // g:/fpga/mxo2/system/project/uart_top.v(84[24:42])
    defparam add_35_5.INIT0 = 16'h5aaa;
    defparam add_35_5.INIT1 = 16'h5aaa;
    defparam add_35_5.INJECT1_0 = "NO";
    defparam add_35_5.INJECT1_1 = "NO";
    CCU2D add_35_3 (.A0(data_length[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(data_length[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n20505), .COUT(n20506), .S0(n78[1]), .S1(n78[2]));   // g:/fpga/mxo2/system/project/uart_top.v(84[24:42])
    defparam add_35_3.INIT0 = 16'h5aaa;
    defparam add_35_3.INIT1 = 16'h5aaa;
    defparam add_35_3.INJECT1_0 = "NO";
    defparam add_35_3.INJECT1_1 = "NO";
    CCU2D add_35_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(data_length[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n20505), .S1(n78[0]));   // g:/fpga/mxo2/system/project/uart_top.v(84[24:42])
    defparam add_35_1.INIT0 = 16'hF000;
    defparam add_35_1.INIT1 = 16'h5555;
    defparam add_35_1.INJECT1_0 = "NO";
    defparam add_35_1.INJECT1_1 = "NO";
    LUT4 i13091_3_lut (.A(tx_data_length[0]), .B(flag), .C(tx_done), .Z(tx_data_length_1__N_1866[0])) /* synthesis lut_function=(A (B+!(C))+!A (B+(C))) */ ;   // g:/fpga/mxo2/system/project/uart_top.v(48[10] 49[49])
    defparam i13091_3_lut.init = 16'hdede;
    LUT4 i2_4_lut (.A(bps_en_tx2), .B(bps_en_tx), .C(bps_en_tx0), .D(bps_en_tx1), 
         .Z(tx_done)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // g:/fpga/mxo2/system/project/uart_top.v(40[18:72])
    defparam i2_4_lut.init = 16'h0200;
    LUT4 i1_2_lut (.A(tx_done), .B(flag), .Z(clk_c_enable_1418)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 tx_data_7__I_0_i1_3_lut (.A(\tamp_data[0] ), .B(\tamp_data[4] ), 
         .C(flag), .Z(tx_data_7__N_1868[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/uart_top.v(58[10] 59[42])
    defparam tx_data_7__I_0_i1_3_lut.init = 16'hcaca;
    LUT4 flag_I_0_4_lut (.A(flag), .B(tx_done), .C(tx_data_length[0]), 
         .D(tx_data_length[1]), .Z(tx_en)) /* synthesis lut_function=(A+(B (C+(D)))) */ ;   // g:/fpga/mxo2/system/project/uart_top.v(63[16:52])
    defparam flag_I_0_4_lut.init = 16'heeea;
    FD1P3IX rx_done_64_rep_506 (.D(n26780), .SP(rx_done_N_2858), .CD(n26803), 
            .CK(clk_c), .Q(n26803)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(101[10] 104[25])
    defparam rx_done_64_rep_506.GSR = "ENABLED";
    FD1P3IX data_length__i1 (.D(n78[1]), .SP(clk_c_enable_1399), .CD(rx_done), 
            .CK(clk_c), .Q(data_length[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(79[10] 84[43])
    defparam data_length__i1.GSR = "ENABLED";
    FD1P3IX data_length__i2 (.D(n78[2]), .SP(clk_c_enable_1399), .CD(rx_done), 
            .CK(clk_c), .Q(data_length[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(79[10] 84[43])
    defparam data_length__i2.GSR = "ENABLED";
    FD1P3IX data_length__i3 (.D(n78[3]), .SP(clk_c_enable_1399), .CD(rx_done), 
            .CK(clk_c), .Q(data_length[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(79[10] 84[43])
    defparam data_length__i3.GSR = "ENABLED";
    FD1P3IX data_length__i4 (.D(n78[4]), .SP(clk_c_enable_1399), .CD(rx_done), 
            .CK(clk_c), .Q(data_length[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(79[10] 84[43])
    defparam data_length__i4.GSR = "ENABLED";
    FD1P3IX data_length__i5 (.D(n78[5]), .SP(clk_c_enable_1399), .CD(rx_done), 
            .CK(clk_c), .Q(data_length[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(79[10] 84[43])
    defparam data_length__i5.GSR = "ENABLED";
    FD1P3IX data_length__i6 (.D(n78[6]), .SP(clk_c_enable_1399), .CD(rx_done), 
            .CK(clk_c), .Q(data_length[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(79[10] 84[43])
    defparam data_length__i6.GSR = "ENABLED";
    FD1P3IX data_length__i7 (.D(n78[7]), .SP(clk_c_enable_1399), .CD(rx_done), 
            .CK(clk_c), .Q(data_length[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(79[10] 84[43])
    defparam data_length__i7.GSR = "ENABLED";
    FD1P3IX data_length__i8 (.D(n78[8]), .SP(clk_c_enable_1399), .CD(rx_done), 
            .CK(clk_c), .Q(data_length[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(79[10] 84[43])
    defparam data_length__i8.GSR = "ENABLED";
    FD1P3IX data_length__i9 (.D(n78[9]), .SP(clk_c_enable_1399), .CD(rx_done), 
            .CK(clk_c), .Q(data_length[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(79[10] 84[43])
    defparam data_length__i9.GSR = "ENABLED";
    FD1P3IX rx_done_64_rep_505 (.D(n26780), .SP(rx_done_N_2858), .CD(n26802), 
            .CK(clk_c), .Q(n26802)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(101[10] 104[25])
    defparam rx_done_64_rep_505.GSR = "ENABLED";
    FD1P3IX rx_done_64_rep_504 (.D(n26780), .SP(rx_done_N_2858), .CD(n26801), 
            .CK(clk_c), .Q(n26801)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(101[10] 104[25])
    defparam rx_done_64_rep_504.GSR = "ENABLED";
    FD1P3IX rx_done_64_rep_503 (.D(n26780), .SP(rx_done_N_2858), .CD(n26800), 
            .CK(clk_c), .Q(n26800)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(101[10] 104[25])
    defparam rx_done_64_rep_503.GSR = "ENABLED";
    LUT4 i1_2_lut_adj_70 (.A(tx_data_length[1]), .B(tx_data_length[0]), 
         .Z(n9394)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i1_2_lut_adj_70.init = 16'h9999;
    LUT4 tx_data_7__I_0_i2_3_lut (.A(\tamp_data[1] ), .B(\tamp_data[5] ), 
         .C(flag), .Z(tx_data_7__N_1868[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/uart_top.v(58[10] 59[42])
    defparam tx_data_7__I_0_i2_3_lut.init = 16'hcaca;
    LUT4 tx_data_7__I_0_i3_3_lut (.A(\tamp_data[2] ), .B(\tamp_data[6] ), 
         .C(flag), .Z(tx_data_7__N_1868[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/uart_top.v(58[10] 59[42])
    defparam tx_data_7__I_0_i3_3_lut.init = 16'hcaca;
    LUT4 tx_data_7__I_0_i4_3_lut (.A(\tamp_data[3] ), .B(\tamp_data[7] ), 
         .C(flag), .Z(tx_data_7__N_1868[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/uart_top.v(58[10] 59[42])
    defparam tx_data_7__I_0_i4_3_lut.init = 16'hcaca;
    FD1P3IX tx_data_i5 (.D(\tamp_data[9] ), .SP(clk_c_enable_1418), .CD(n12084), 
            .CK(clk_c), .Q(tx_data[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(56[10] 59[42])
    defparam tx_data_i5.GSR = "ENABLED";
    FD1P3IX tx_data_i4 (.D(\tamp_data[8] ), .SP(clk_c_enable_1418), .CD(n12084), 
            .CK(clk_c), .Q(tx_data[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(56[10] 59[42])
    defparam tx_data_i4.GSR = "ENABLED";
    LUT4 i7_4_lut (.A(n9), .B(n23801), .C(rx_data[5]), .D(rx_data[2]), 
         .Z(n15)) /* synthesis lut_function=(A+((C+!(D))+!B)) */ ;
    defparam i7_4_lut.init = 16'hfbff;
    LUT4 i1_2_lut_adj_71 (.A(rx_data[6]), .B(rx_data[7]), .Z(n9)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_71.init = 16'heeee;
    LUT4 i20925_4_lut (.A(rx_data[3]), .B(rx_data[0]), .C(rx_data[1]), 
         .D(rx_data[4]), .Z(n23801)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i20925_4_lut.init = 16'h8000;
    FD1P3IX rx_done_64_rep_502 (.D(n26780), .SP(rx_done_N_2858), .CD(n26799), 
            .CK(clk_c), .Q(n26799)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(101[10] 104[25])
    defparam rx_done_64_rep_502.GSR = "ENABLED";
    LUT4 ready_I_0_2_lut (.A(ready), .B(n15), .Z(rx_done_N_2858)) /* synthesis lut_function=(!((B)+!A)) */ ;   // g:/fpga/mxo2/system/project/uart_top.v(81[15:38])
    defparam ready_I_0_2_lut.init = 16'h2222;
    FD1P3IX rx_done_64_rep_501 (.D(n26780), .SP(rx_done_N_2858), .CD(n26798), 
            .CK(clk_c), .Q(n26798)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(101[10] 104[25])
    defparam rx_done_64_rep_501.GSR = "ENABLED";
    FD1P3IX rx_done_64_rep_500 (.D(n26780), .SP(rx_done_N_2858), .CD(n26797), 
            .CK(clk_c), .Q(n26797)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(101[10] 104[25])
    defparam rx_done_64_rep_500.GSR = "ENABLED";
    FD1P3IX rx_done_64_rep_499 (.D(n26780), .SP(rx_done_N_2858), .CD(n26796), 
            .CK(clk_c), .Q(n26796)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(101[10] 104[25])
    defparam rx_done_64_rep_499.GSR = "ENABLED";
    FD1P3IX rx_done_64_rep_498 (.D(n26780), .SP(rx_done_N_2858), .CD(n26795), 
            .CK(clk_c), .Q(n26795)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=91, LSE_RLINE=101 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(101[10] 104[25])
    defparam rx_done_64_rep_498.GSR = "ENABLED";
    uart_tx uart_tx_ins (.clk_c(clk_c), .bps_en_N_2978(bps_en_N_2978), .\tx_data[0] (tx_data[0]), 
            .bps_en_tx(bps_en_tx), .bps_clk_tx(bps_clk_tx), .rs232_tx_c(rs232_tx_c), 
            .\tx_data[1] (tx_data[1]), .\tx_data[2] (tx_data[2]), .\tx_data[3] (tx_data[3]), 
            .\tx_data[4] (tx_data[4]), .\tx_data[5] (tx_data[5]), .n26780(n26780)) /* synthesis syn_module_defined=1 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(150[9] 159[2])
    uart_rx uart_rx_ins (.rx_data({rx_data}), .clk_c(clk_c), .bps_en_rx(bps_en_rx), 
            .rs232_rx_c(rs232_rx_c), .ready(ready), .n26780(n26780), .bps_clk_rx(bps_clk_rx)) /* synthesis syn_module_defined=1 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(123[9] 132[2])
    baud_generator baud_tx_ins (.bps_clk_tx(bps_clk_tx), .clk_c(clk_c), 
            .GND_net(GND_net), .bps_en_tx(bps_en_tx)) /* synthesis syn_module_defined=1 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(141[1] 147[2])
    baud_generator_U0 baud_rx_ins (.bps_clk_rx(bps_clk_rx), .clk_c(clk_c), 
            .bps_en_rx(bps_en_rx), .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // g:/fpga/mxo2/system/project/uart_top.v(114[1] 120[2])
    
endmodule
//
// Verilog Description of module uart_tx
//

module uart_tx (clk_c, bps_en_N_2978, \tx_data[0] , bps_en_tx, bps_clk_tx, 
            rs232_tx_c, \tx_data[1] , \tx_data[2] , \tx_data[3] , \tx_data[4] , 
            \tx_data[5] , n26780) /* synthesis syn_module_defined=1 */ ;
    input clk_c;
    input bps_en_N_2978;
    input \tx_data[0] ;
    output bps_en_tx;
    input bps_clk_tx;
    output rs232_tx_c;
    input \tx_data[1] ;
    input \tx_data[2] ;
    input \tx_data[3] ;
    input \tx_data[4] ;
    input \tx_data[5] ;
    input n26780;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // g:/fpga/mxo2/system/project/system_top.v(2[15:18])
    wire [3:0]num;   // g:/fpga/mxo2/system/project/uart_tx.v(12[14:17])
    
    wire n8719;
    wire [10:0]tx_data_r;   // g:/fpga/mxo2/system/project/uart_tx.v(13[15:24])
    
    wire n11846, clk_c_enable_1358, n12038, n1, n7, n24611, clk_c_enable_687, 
        rs232_tx_N_2983;
    wire [3:0]n21;
    
    wire n24612, n24613, n24615, n2, n1_adj_5031, n23882, n24614;
    
    LUT4 i6129_2_lut (.A(num[0]), .B(num[1]), .Z(n8719)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // g:/fpga/mxo2/system/project/uart_tx.v(35[26:29])
    defparam i6129_2_lut.init = 16'h6666;
    FD1P3AX tx_data_r__i1 (.D(\tx_data[0] ), .SP(bps_en_N_2978), .CK(clk_c), 
            .Q(tx_data_r[1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=150, LSE_RLINE=159 */ ;   // g:/fpga/mxo2/system/project/uart_tx.v(19[11] 24[5])
    defparam tx_data_r__i1.GSR = "ENABLED";
    FD1S3AX bps_en_24 (.D(n11846), .CK(clk_c), .Q(bps_en_tx)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=150, LSE_RLINE=159 */ ;   // g:/fpga/mxo2/system/project/uart_tx.v(19[11] 24[5])
    defparam bps_en_24.GSR = "ENABLED";
    FD1P3IX num_1986__i0 (.D(n1), .SP(clk_c_enable_1358), .CD(n12038), 
            .CK(clk_c), .Q(num[0]));   // g:/fpga/mxo2/system/project/uart_tx.v(34[11:21])
    defparam num_1986__i0.GSR = "ENABLED";
    LUT4 i21577_3_lut_rep_372 (.A(n7), .B(bps_en_tx), .C(bps_clk_tx), 
         .Z(clk_c_enable_1358)) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;
    defparam i21577_3_lut_rep_372.init = 16'hc4c4;
    LUT4 i21445_2_lut_3_lut (.A(n7), .B(bps_en_tx), .C(bps_clk_tx), .Z(n12038)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;
    defparam i21445_2_lut_3_lut.init = 16'h0404;
    LUT4 n23882_bdd_4_lut_22120 (.A(num[0]), .B(num[1]), .C(tx_data_r[10]), 
         .D(num[2]), .Z(n24611)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (((D)+!C)+!B))) */ ;
    defparam n23882_bdd_4_lut_22120.init = 16'h0060;
    FD1P3AY rs232_tx_28 (.D(rs232_tx_N_2983), .SP(clk_c_enable_687), .CK(clk_c), 
            .Q(rs232_tx_c)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=150, LSE_RLINE=159 */ ;   // g:/fpga/mxo2/system/project/uart_tx.v(32[11] 38[5])
    defparam rs232_tx_28.GSR = "ENABLED";
    FD1P3IX num_1986__i3 (.D(n21[3]), .SP(clk_c_enable_1358), .CD(n12038), 
            .CK(clk_c), .Q(num[3]));   // g:/fpga/mxo2/system/project/uart_tx.v(34[11:21])
    defparam num_1986__i3.GSR = "ENABLED";
    FD1P3IX num_1986__i2 (.D(n21[2]), .SP(clk_c_enable_1358), .CD(n12038), 
            .CK(clk_c), .Q(num[2]));   // g:/fpga/mxo2/system/project/uart_tx.v(34[11:21])
    defparam num_1986__i2.GSR = "ENABLED";
    FD1P3IX num_1986__i1 (.D(n8719), .SP(clk_c_enable_1358), .CD(n12038), 
            .CK(clk_c), .Q(num[1]));   // g:/fpga/mxo2/system/project/uart_tx.v(34[11:21])
    defparam num_1986__i1.GSR = "ENABLED";
    LUT4 i17642_3_lut_4_lut (.A(num[1]), .B(num[0]), .C(num[2]), .D(num[3]), 
         .Z(n21[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // g:/fpga/mxo2/system/project/uart_tx.v(34[11:21])
    defparam i17642_3_lut_4_lut.init = 16'h7f80;
    FD1P3AX tx_data_r__i2 (.D(\tx_data[1] ), .SP(bps_en_N_2978), .CK(clk_c), 
            .Q(tx_data_r[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=150, LSE_RLINE=159 */ ;   // g:/fpga/mxo2/system/project/uart_tx.v(19[11] 24[5])
    defparam tx_data_r__i2.GSR = "ENABLED";
    FD1P3AX tx_data_r__i3 (.D(\tx_data[2] ), .SP(bps_en_N_2978), .CK(clk_c), 
            .Q(tx_data_r[3])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=150, LSE_RLINE=159 */ ;   // g:/fpga/mxo2/system/project/uart_tx.v(19[11] 24[5])
    defparam tx_data_r__i3.GSR = "ENABLED";
    FD1P3AX tx_data_r__i4 (.D(\tx_data[3] ), .SP(bps_en_N_2978), .CK(clk_c), 
            .Q(tx_data_r[4])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=150, LSE_RLINE=159 */ ;   // g:/fpga/mxo2/system/project/uart_tx.v(19[11] 24[5])
    defparam tx_data_r__i4.GSR = "ENABLED";
    FD1P3AX tx_data_r__i5 (.D(\tx_data[4] ), .SP(bps_en_N_2978), .CK(clk_c), 
            .Q(tx_data_r[5])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=150, LSE_RLINE=159 */ ;   // g:/fpga/mxo2/system/project/uart_tx.v(19[11] 24[5])
    defparam tx_data_r__i5.GSR = "ENABLED";
    FD1P3AX tx_data_r__i6 (.D(\tx_data[5] ), .SP(bps_en_N_2978), .CK(clk_c), 
            .Q(tx_data_r[6])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=150, LSE_RLINE=159 */ ;   // g:/fpga/mxo2/system/project/uart_tx.v(19[11] 24[5])
    defparam tx_data_r__i6.GSR = "ENABLED";
    FD1P3AX tx_data_r__i9 (.D(n26780), .SP(bps_en_N_2978), .CK(clk_c), 
            .Q(tx_data_r[10])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=150, LSE_RLINE=159 */ ;   // g:/fpga/mxo2/system/project/uart_tx.v(19[11] 24[5])
    defparam tx_data_r__i9.GSR = "ENABLED";
    LUT4 i9035_3_lut (.A(n7), .B(bps_en_N_2978), .C(bps_en_tx), .Z(n11846)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;   // g:/fpga/mxo2/system/project/uart_tx.v(19[11] 24[5])
    defparam i9035_3_lut.init = 16'hecec;
    LUT4 i2_4_lut (.A(num[3]), .B(num[2]), .C(num[1]), .D(num[0]), .Z(n7)) /* synthesis lut_function=((B+!(C (D)))+!A) */ ;
    defparam i2_4_lut.init = 16'hdfff;
    LUT4 i2908_1_lut (.A(num[0]), .Z(n1)) /* synthesis lut_function=(!(A)) */ ;   // g:/fpga/mxo2/system/project/uart_tx.v(22[14:24])
    defparam i2908_1_lut.init = 16'h5555;
    LUT4 i17635_2_lut_3_lut (.A(num[1]), .B(num[0]), .C(num[2]), .Z(n21[2])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // g:/fpga/mxo2/system/project/uart_tx.v(34[11:21])
    defparam i17635_2_lut_3_lut.init = 16'h7878;
    LUT4 tx_data_r_5__bdd_2_lut_22121 (.A(tx_data_r[5]), .B(num[1]), .Z(n24612)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam tx_data_r_5__bdd_2_lut_22121.init = 16'h2222;
    LUT4 tx_data_r_5__bdd_3_lut_22122 (.A(tx_data_r[4]), .B(num[1]), .C(tx_data_r[6]), 
         .Z(n24613)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam tx_data_r_5__bdd_3_lut_22122.init = 16'he2e2;
    LUT4 i3157_2_lut (.A(bps_clk_tx), .B(bps_en_tx), .Z(clk_c_enable_687)) /* synthesis lut_function=(A (B)) */ ;   // g:/fpga/mxo2/system/project/uart_tx.v(32[11] 38[5])
    defparam i3157_2_lut.init = 16'h8888;
    LUT4 n24615_bdd_3_lut (.A(n24615), .B(n24611), .C(num[3]), .Z(rs232_tx_N_2983)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24615_bdd_3_lut.init = 16'hcaca;
    LUT4 num_3__I_0_i2_3_lut (.A(tx_data_r[2]), .B(tx_data_r[3]), .C(num[0]), 
         .Z(n2)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/uart_tx.v(35[26:29])
    defparam num_3__I_0_i2_3_lut.init = 16'hcaca;
    LUT4 i13096_2_lut (.A(tx_data_r[1]), .B(num[0]), .Z(n1_adj_5031)) /* synthesis lut_function=(A (B)) */ ;   // g:/fpga/mxo2/system/project/uart_tx.v(35[26:29])
    defparam i13096_2_lut.init = 16'h8888;
    PFUMX i21005 (.BLUT(n1_adj_5031), .ALUT(n2), .C0(num[1]), .Z(n23882));
    L6MUX21 i21619 (.D0(n23882), .D1(n24614), .SD(num[2]), .Z(n24615));
    PFUMX i21617 (.BLUT(n24613), .ALUT(n24612), .C0(num[0]), .Z(n24614));
    
endmodule
//
// Verilog Description of module uart_rx
//

module uart_rx (rx_data, clk_c, bps_en_rx, rs232_rx_c, ready, n26780, 
            bps_clk_rx) /* synthesis syn_module_defined=1 */ ;
    output [7:0]rx_data;
    input clk_c;
    output bps_en_rx;
    input rs232_rx_c;
    output ready;
    input n26780;
    input bps_clk_rx;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // g:/fpga/mxo2/system/project/system_top.v(2[15:18])
    
    wire clk_c_enable_743;
    wire [7:0]rx_data_r;   // g:/fpga/mxo2/system/project/uart_rx.v(42[14:23])
    
    wire rs232_rx1, rs232_rx0, rs232_rx2, n11848;
    wire [3:0]num;   // g:/fpga/mxo2/system/project/uart_rx.v(31[14:17])
    
    wire clk_c_enable_1362, n12037;
    wire [3:0]n21;
    
    wire bps_en_N_2945, n9142, clk_c_enable_1404, clk_c_enable_1406, 
        clk_c_enable_1405, clk_c_enable_1403, n16586, n23227, clk_c_enable_1379, 
        clk_c_enable_1402, clk_c_enable_1407, clk_c_enable_1408;
    
    FD1P3AX rx_data_i0_i0 (.D(rx_data_r[0]), .SP(clk_c_enable_743), .CK(clk_c), 
            .Q(rx_data[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=132 */ ;   // g:/fpga/mxo2/system/project/uart_rx.v(49[11] 58[5])
    defparam rx_data_i0_i0.GSR = "ENABLED";
    FD1S3AX rs232_rx1_56 (.D(rs232_rx0), .CK(clk_c), .Q(rs232_rx1)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=132 */ ;   // g:/fpga/mxo2/system/project/uart_rx.v(21[11] 25[5])
    defparam rs232_rx1_56.GSR = "ENABLED";
    FD1S3AX rs232_rx2_57 (.D(rs232_rx1), .CK(clk_c), .Q(rs232_rx2)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=132 */ ;   // g:/fpga/mxo2/system/project/uart_rx.v(21[11] 25[5])
    defparam rs232_rx2_57.GSR = "ENABLED";
    FD1S3AX bps_en_58 (.D(n11848), .CK(clk_c), .Q(bps_en_rx)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=132 */ ;   // g:/fpga/mxo2/system/project/uart_rx.v(36[7] 39[18])
    defparam bps_en_58.GSR = "ENABLED";
    FD1S3AX rs232_rx0_55 (.D(rs232_rx_c), .CK(clk_c), .Q(rs232_rx0)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=132 */ ;   // g:/fpga/mxo2/system/project/uart_rx.v(21[11] 25[5])
    defparam rs232_rx0_55.GSR = "ENABLED";
    FD1P3IX num_1984__i0 (.D(n21[0]), .SP(clk_c_enable_1362), .CD(n12037), 
            .CK(clk_c), .Q(num[0]));   // g:/fpga/mxo2/system/project/uart_rx.v(51[11:19])
    defparam num_1984__i0.GSR = "ENABLED";
    FD1P3IX ready_62 (.D(n26780), .SP(bps_en_N_2945), .CD(ready), .CK(clk_c), 
            .Q(ready)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=132 */ ;   // g:/fpga/mxo2/system/project/uart_rx.v(64[10] 67[23])
    defparam ready_62.GSR = "ENABLED";
    LUT4 i21532_2_lut_3_lut_4_lut (.A(n9142), .B(num[0]), .C(num[1]), 
         .D(num[2]), .Z(clk_c_enable_1404)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // g:/fpga/mxo2/system/project/uart_rx.v(53[4:20])
    defparam i21532_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i17599_2_lut (.A(num[1]), .B(num[0]), .Z(n21[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // g:/fpga/mxo2/system/project/uart_rx.v(51[11:19])
    defparam i17599_2_lut.init = 16'h6666;
    LUT4 i21528_2_lut_3_lut_4_lut (.A(n9142), .B(num[0]), .C(num[1]), 
         .D(num[2]), .Z(clk_c_enable_1406)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // g:/fpga/mxo2/system/project/uart_rx.v(53[4:20])
    defparam i21528_2_lut_3_lut_4_lut.init = 16'h0200;
    LUT4 i21530_2_lut_3_lut_4_lut (.A(n9142), .B(num[0]), .C(num[1]), 
         .D(num[2]), .Z(clk_c_enable_1405)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i21530_2_lut_3_lut_4_lut.init = 16'h0800;
    LUT4 i13942_2_lut_3_lut_4_lut (.A(n9142), .B(num[0]), .C(num[1]), 
         .D(num[2]), .Z(clk_c_enable_1403)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i13942_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i2_3_lut (.A(bps_en_rx), .B(bps_clk_rx), .C(bps_en_N_2945), .Z(clk_c_enable_743)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // g:/fpga/mxo2/system/project/uart_rx.v(49[11] 58[5])
    defparam i2_3_lut.init = 16'h2020;
    LUT4 i2_4_lut (.A(bps_en_rx), .B(bps_clk_rx), .C(n16586), .D(num[3]), 
         .Z(n9142)) /* synthesis lut_function=(!(((C (D))+!B)+!A)) */ ;   // g:/fpga/mxo2/system/project/uart_rx.v(49[11] 58[5])
    defparam i2_4_lut.init = 16'h0888;
    FD1P3AX rx_data_i0_i1 (.D(rx_data_r[1]), .SP(clk_c_enable_743), .CK(clk_c), 
            .Q(rx_data[1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=132 */ ;   // g:/fpga/mxo2/system/project/uart_rx.v(49[11] 58[5])
    defparam rx_data_i0_i1.GSR = "ENABLED";
    FD1P3AX rx_data_i0_i2 (.D(rx_data_r[2]), .SP(clk_c_enable_743), .CK(clk_c), 
            .Q(rx_data[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=132 */ ;   // g:/fpga/mxo2/system/project/uart_rx.v(49[11] 58[5])
    defparam rx_data_i0_i2.GSR = "ENABLED";
    FD1P3AX rx_data_i0_i3 (.D(rx_data_r[3]), .SP(clk_c_enable_743), .CK(clk_c), 
            .Q(rx_data[3])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=132 */ ;   // g:/fpga/mxo2/system/project/uart_rx.v(49[11] 58[5])
    defparam rx_data_i0_i3.GSR = "ENABLED";
    FD1P3AX rx_data_i0_i4 (.D(rx_data_r[4]), .SP(clk_c_enable_743), .CK(clk_c), 
            .Q(rx_data[4])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=132 */ ;   // g:/fpga/mxo2/system/project/uart_rx.v(49[11] 58[5])
    defparam rx_data_i0_i4.GSR = "ENABLED";
    FD1P3AX rx_data_i0_i5 (.D(rx_data_r[5]), .SP(clk_c_enable_743), .CK(clk_c), 
            .Q(rx_data[5])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=132 */ ;   // g:/fpga/mxo2/system/project/uart_rx.v(49[11] 58[5])
    defparam rx_data_i0_i5.GSR = "ENABLED";
    FD1P3AX rx_data_i0_i6 (.D(rx_data_r[6]), .SP(clk_c_enable_743), .CK(clk_c), 
            .Q(rx_data[6])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=132 */ ;   // g:/fpga/mxo2/system/project/uart_rx.v(49[11] 58[5])
    defparam rx_data_i0_i6.GSR = "ENABLED";
    FD1P3AX rx_data_i0_i7 (.D(rx_data_r[7]), .SP(clk_c_enable_743), .CK(clk_c), 
            .Q(rx_data[7])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=132 */ ;   // g:/fpga/mxo2/system/project/uart_rx.v(49[11] 58[5])
    defparam rx_data_i0_i7.GSR = "ENABLED";
    LUT4 i21580_3_lut_rep_329 (.A(bps_en_N_2945), .B(bps_en_rx), .C(bps_clk_rx), 
         .Z(clk_c_enable_1362)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i21580_3_lut_rep_329.init = 16'hc8c8;
    LUT4 i21439_2_lut_3_lut (.A(bps_en_N_2945), .B(bps_en_rx), .C(bps_clk_rx), 
         .Z(n12037)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i21439_2_lut_3_lut.init = 16'h0808;
    FD1P3IX num_1984__i3 (.D(n21[3]), .SP(clk_c_enable_1362), .CD(n12037), 
            .CK(clk_c), .Q(num[3]));   // g:/fpga/mxo2/system/project/uart_rx.v(51[11:19])
    defparam num_1984__i3.GSR = "ENABLED";
    FD1P3IX num_1984__i2 (.D(n21[2]), .SP(clk_c_enable_1362), .CD(n12037), 
            .CK(clk_c), .Q(num[2]));   // g:/fpga/mxo2/system/project/uart_rx.v(51[11:19])
    defparam num_1984__i2.GSR = "ENABLED";
    FD1P3IX num_1984__i1 (.D(n21[1]), .SP(clk_c_enable_1362), .CD(n12037), 
            .CK(clk_c), .Q(num[1]));   // g:/fpga/mxo2/system/project/uart_rx.v(51[11:19])
    defparam num_1984__i1.GSR = "ENABLED";
    LUT4 i9037_4_lut (.A(bps_en_N_2945), .B(n23227), .C(bps_en_rx), .D(rs232_rx1), 
         .Z(n11848)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A !(B (C+(D))+!B (C)))) */ ;   // g:/fpga/mxo2/system/project/uart_rx.v(36[7] 39[18])
    defparam i9037_4_lut.init = 16'h5c50;
    LUT4 i2_3_lut_adj_69 (.A(rs232_rx_c), .B(rs232_rx0), .C(rs232_rx2), 
         .Z(n23227)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // g:/fpga/mxo2/system/project/uart_rx.v(36[10:35])
    defparam i2_3_lut_adj_69.init = 16'h1010;
    LUT4 i21458_3_lut_4_lut (.A(num[1]), .B(num[2]), .C(num[0]), .D(num[3]), 
         .Z(bps_en_N_2945)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // g:/fpga/mxo2/system/project/uart_rx.v(53[4:20])
    defparam i21458_3_lut_4_lut.init = 16'h1000;
    LUT4 i13801_2_lut_3_lut (.A(num[1]), .B(num[2]), .C(num[0]), .Z(n16586)) /* synthesis lut_function=(A+(B+(C))) */ ;   // g:/fpga/mxo2/system/project/uart_rx.v(53[4:20])
    defparam i13801_2_lut_3_lut.init = 16'hfefe;
    LUT4 i21343_2_lut_3_lut_3_lut_4_lut (.A(num[1]), .B(num[2]), .C(n9142), 
         .D(num[0]), .Z(clk_c_enable_1379)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // g:/fpga/mxo2/system/project/uart_rx.v(53[4:20])
    defparam i21343_2_lut_3_lut_3_lut_4_lut.init = 16'h1000;
    FD1P3AX rx_data_r_i0_i0 (.D(rs232_rx_c), .SP(clk_c_enable_1379), .CK(clk_c), 
            .Q(rx_data_r[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=132 */ ;   // g:/fpga/mxo2/system/project/uart_rx.v(49[11] 58[5])
    defparam rx_data_r_i0_i0.GSR = "ENABLED";
    LUT4 i21535_2_lut_2_lut_3_lut_4_lut (.A(num[1]), .B(num[2]), .C(num[0]), 
         .D(n9142), .Z(clk_c_enable_1402)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // g:/fpga/mxo2/system/project/uart_rx.v(53[4:20])
    defparam i21535_2_lut_2_lut_3_lut_4_lut.init = 16'h0100;
    FD1P3AX rx_data_r_i0_i7 (.D(rs232_rx_c), .SP(clk_c_enable_1402), .CK(clk_c), 
            .Q(rx_data_r[7])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=132 */ ;   // g:/fpga/mxo2/system/project/uart_rx.v(49[11] 58[5])
    defparam rx_data_r_i0_i7.GSR = "ENABLED";
    FD1P3AX rx_data_r_i0_i6 (.D(rs232_rx_c), .SP(clk_c_enable_1403), .CK(clk_c), 
            .Q(rx_data_r[6])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=132 */ ;   // g:/fpga/mxo2/system/project/uart_rx.v(49[11] 58[5])
    defparam rx_data_r_i0_i6.GSR = "ENABLED";
    FD1P3AX rx_data_r_i0_i5 (.D(rs232_rx_c), .SP(clk_c_enable_1404), .CK(clk_c), 
            .Q(rx_data_r[5])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=132 */ ;   // g:/fpga/mxo2/system/project/uart_rx.v(49[11] 58[5])
    defparam rx_data_r_i0_i5.GSR = "ENABLED";
    FD1P3AX rx_data_r_i0_i4 (.D(rs232_rx_c), .SP(clk_c_enable_1405), .CK(clk_c), 
            .Q(rx_data_r[4])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=132 */ ;   // g:/fpga/mxo2/system/project/uart_rx.v(49[11] 58[5])
    defparam rx_data_r_i0_i4.GSR = "ENABLED";
    FD1P3AX rx_data_r_i0_i3 (.D(rs232_rx_c), .SP(clk_c_enable_1406), .CK(clk_c), 
            .Q(rx_data_r[3])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=132 */ ;   // g:/fpga/mxo2/system/project/uart_rx.v(49[11] 58[5])
    defparam rx_data_r_i0_i3.GSR = "ENABLED";
    FD1P3AX rx_data_r_i0_i2 (.D(rs232_rx_c), .SP(clk_c_enable_1407), .CK(clk_c), 
            .Q(rx_data_r[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=132 */ ;   // g:/fpga/mxo2/system/project/uart_rx.v(49[11] 58[5])
    defparam rx_data_r_i0_i2.GSR = "ENABLED";
    FD1P3AX rx_data_r_i0_i1 (.D(rs232_rx_c), .SP(clk_c_enable_1408), .CK(clk_c), 
            .Q(rx_data_r[1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=132 */ ;   // g:/fpga/mxo2/system/project/uart_rx.v(49[11] 58[5])
    defparam rx_data_r_i0_i1.GSR = "ENABLED";
    LUT4 i17597_1_lut (.A(num[0]), .Z(n21[0])) /* synthesis lut_function=(!(A)) */ ;   // g:/fpga/mxo2/system/project/uart_rx.v(51[11:19])
    defparam i17597_1_lut.init = 16'h5555;
    LUT4 i21496_2_lut_3_lut_3_lut_4_lut (.A(num[2]), .B(num[1]), .C(n9142), 
         .D(num[0]), .Z(clk_c_enable_1408)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // g:/fpga/mxo2/system/project/uart_rx.v(53[4:20])
    defparam i21496_2_lut_3_lut_3_lut_4_lut.init = 16'h0040;
    LUT4 i21525_2_lut_3_lut_3_lut_4_lut (.A(num[2]), .B(num[1]), .C(n9142), 
         .D(num[0]), .Z(clk_c_enable_1407)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // g:/fpga/mxo2/system/project/uart_rx.v(53[4:20])
    defparam i21525_2_lut_3_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 i17613_3_lut_4_lut (.A(num[1]), .B(num[0]), .C(num[2]), .D(num[3]), 
         .Z(n21[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // g:/fpga/mxo2/system/project/uart_rx.v(51[11:19])
    defparam i17613_3_lut_4_lut.init = 16'h7f80;
    LUT4 i17606_2_lut_3_lut (.A(num[1]), .B(num[0]), .C(num[2]), .Z(n21[2])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // g:/fpga/mxo2/system/project/uart_rx.v(51[11:19])
    defparam i17606_2_lut_3_lut.init = 16'h7878;
    
endmodule
//
// Verilog Description of module baud_generator
//

module baud_generator (bps_clk_tx, clk_c, GND_net, bps_en_tx) /* synthesis syn_module_defined=1 */ ;
    output bps_clk_tx;
    input clk_c;
    input GND_net;
    input bps_en_tx;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // g:/fpga/mxo2/system/project/system_top.v(2[15:18])
    
    wire bps_clk_N_2900;
    wire [12:0]cnt;   // g:/fpga/mxo2/system/project/baud_generator.v(12[15:18])
    
    wire cnt_12__N_2896;
    wire [12:0]n57;
    
    wire n25732, n7, n23618, n8, n23123, n20560, n20559, n20558, 
        n20853, n5, n6, n20557, n20556, n20555;
    
    FD1S3AX bps_clk_17 (.D(bps_clk_N_2900), .CK(clk_c), .Q(bps_clk_tx)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=141, LSE_RLINE=147 */ ;   // g:/fpga/mxo2/system/project/baud_generator.v(28[8] 31[20])
    defparam bps_clk_17.GSR = "ENABLED";
    FD1S3IX cnt_1985__i0 (.D(n57[0]), .CK(clk_c), .CD(cnt_12__N_2896), 
            .Q(cnt[0])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/baud_generator.v(20[10:20])
    defparam cnt_1985__i0.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_450 (.A(cnt[12]), .B(cnt[11]), .Z(n25732)) /* synthesis lut_function=(A+(B)) */ ;   // g:/fpga/mxo2/system/project/baud_generator.v(17[10:40])
    defparam i1_2_lut_rep_450.init = 16'heeee;
    LUT4 i21453_4_lut (.A(cnt[0]), .B(n7), .C(cnt[6]), .D(n23618), .Z(bps_clk_N_2900)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // g:/fpga/mxo2/system/project/baud_generator.v(28[11:31])
    defparam i21453_4_lut.init = 16'h2000;
    LUT4 i3_3_lut_4_lut (.A(cnt[12]), .B(cnt[11]), .C(cnt[10]), .D(cnt[7]), 
         .Z(n8)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // g:/fpga/mxo2/system/project/baud_generator.v(17[10:40])
    defparam i3_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut (.A(cnt[9]), .B(cnt[8]), .C(n8), .D(n23123), .Z(n7)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i1_4_lut.init = 16'hfffd;
    LUT4 i20759_2_lut (.A(cnt[5]), .B(cnt[4]), .Z(n23618)) /* synthesis lut_function=(A (B)) */ ;
    defparam i20759_2_lut.init = 16'h8888;
    LUT4 i2_3_lut (.A(cnt[1]), .B(cnt[2]), .C(cnt[3]), .Z(n23123)) /* synthesis lut_function=(A+(B+(C))) */ ;   // g:/fpga/mxo2/system/project/baud_generator.v(17[10:40])
    defparam i2_3_lut.init = 16'hfefe;
    FD1S3IX cnt_1985__i1 (.D(n57[1]), .CK(clk_c), .CD(cnt_12__N_2896), 
            .Q(cnt[1])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/baud_generator.v(20[10:20])
    defparam cnt_1985__i1.GSR = "ENABLED";
    FD1S3IX cnt_1985__i2 (.D(n57[2]), .CK(clk_c), .CD(cnt_12__N_2896), 
            .Q(cnt[2])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/baud_generator.v(20[10:20])
    defparam cnt_1985__i2.GSR = "ENABLED";
    FD1S3IX cnt_1985__i3 (.D(n57[3]), .CK(clk_c), .CD(cnt_12__N_2896), 
            .Q(cnt[3])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/baud_generator.v(20[10:20])
    defparam cnt_1985__i3.GSR = "ENABLED";
    FD1S3IX cnt_1985__i4 (.D(n57[4]), .CK(clk_c), .CD(cnt_12__N_2896), 
            .Q(cnt[4])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/baud_generator.v(20[10:20])
    defparam cnt_1985__i4.GSR = "ENABLED";
    FD1S3IX cnt_1985__i5 (.D(n57[5]), .CK(clk_c), .CD(cnt_12__N_2896), 
            .Q(cnt[5])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/baud_generator.v(20[10:20])
    defparam cnt_1985__i5.GSR = "ENABLED";
    FD1S3IX cnt_1985__i6 (.D(n57[6]), .CK(clk_c), .CD(cnt_12__N_2896), 
            .Q(cnt[6])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/baud_generator.v(20[10:20])
    defparam cnt_1985__i6.GSR = "ENABLED";
    FD1S3IX cnt_1985__i7 (.D(n57[7]), .CK(clk_c), .CD(cnt_12__N_2896), 
            .Q(cnt[7])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/baud_generator.v(20[10:20])
    defparam cnt_1985__i7.GSR = "ENABLED";
    FD1S3IX cnt_1985__i8 (.D(n57[8]), .CK(clk_c), .CD(cnt_12__N_2896), 
            .Q(cnt[8])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/baud_generator.v(20[10:20])
    defparam cnt_1985__i8.GSR = "ENABLED";
    FD1S3IX cnt_1985__i9 (.D(n57[9]), .CK(clk_c), .CD(cnt_12__N_2896), 
            .Q(cnt[9])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/baud_generator.v(20[10:20])
    defparam cnt_1985__i9.GSR = "ENABLED";
    FD1S3IX cnt_1985__i10 (.D(n57[10]), .CK(clk_c), .CD(cnt_12__N_2896), 
            .Q(cnt[10])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/baud_generator.v(20[10:20])
    defparam cnt_1985__i10.GSR = "ENABLED";
    FD1S3IX cnt_1985__i11 (.D(n57[11]), .CK(clk_c), .CD(cnt_12__N_2896), 
            .Q(cnt[11])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/baud_generator.v(20[10:20])
    defparam cnt_1985__i11.GSR = "ENABLED";
    FD1S3IX cnt_1985__i12 (.D(n57[12]), .CK(clk_c), .CD(cnt_12__N_2896), 
            .Q(cnt[12])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/baud_generator.v(20[10:20])
    defparam cnt_1985__i12.GSR = "ENABLED";
    CCU2D cnt_1985_add_4_13 (.A0(cnt[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n20560), .S0(n57[11]), .S1(n57[12]));   // g:/fpga/mxo2/system/project/baud_generator.v(20[10:20])
    defparam cnt_1985_add_4_13.INIT0 = 16'hfaaa;
    defparam cnt_1985_add_4_13.INIT1 = 16'hfaaa;
    defparam cnt_1985_add_4_13.INJECT1_0 = "NO";
    defparam cnt_1985_add_4_13.INJECT1_1 = "NO";
    CCU2D cnt_1985_add_4_11 (.A0(cnt[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n20559), .COUT(n20560), .S0(n57[9]), .S1(n57[10]));   // g:/fpga/mxo2/system/project/baud_generator.v(20[10:20])
    defparam cnt_1985_add_4_11.INIT0 = 16'hfaaa;
    defparam cnt_1985_add_4_11.INIT1 = 16'hfaaa;
    defparam cnt_1985_add_4_11.INJECT1_0 = "NO";
    defparam cnt_1985_add_4_11.INJECT1_1 = "NO";
    CCU2D cnt_1985_add_4_9 (.A0(cnt[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n20558), 
          .COUT(n20559), .S0(n57[7]), .S1(n57[8]));   // g:/fpga/mxo2/system/project/baud_generator.v(20[10:20])
    defparam cnt_1985_add_4_9.INIT0 = 16'hfaaa;
    defparam cnt_1985_add_4_9.INIT1 = 16'hfaaa;
    defparam cnt_1985_add_4_9.INJECT1_0 = "NO";
    defparam cnt_1985_add_4_9.INJECT1_1 = "NO";
    LUT4 i2_4_lut (.A(n25732), .B(n20853), .C(bps_en_tx), .D(cnt[10]), 
         .Z(cnt_12__N_2896)) /* synthesis lut_function=(A+(B ((D)+!C)+!B !(C))) */ ;   // g:/fpga/mxo2/system/project/baud_generator.v(17[10:40])
    defparam i2_4_lut.init = 16'hefaf;
    LUT4 i2_4_lut_adj_67 (.A(cnt[9]), .B(cnt[8]), .C(n5), .D(n6), .Z(n20853)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_67.init = 16'hfeee;
    CCU2D cnt_1985_add_4_7 (.A0(cnt[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n20557), 
          .COUT(n20558), .S0(n57[5]), .S1(n57[6]));   // g:/fpga/mxo2/system/project/baud_generator.v(20[10:20])
    defparam cnt_1985_add_4_7.INIT0 = 16'hfaaa;
    defparam cnt_1985_add_4_7.INIT1 = 16'hfaaa;
    defparam cnt_1985_add_4_7.INJECT1_0 = "NO";
    defparam cnt_1985_add_4_7.INJECT1_1 = "NO";
    CCU2D cnt_1985_add_4_5 (.A0(cnt[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n20556), 
          .COUT(n20557), .S0(n57[3]), .S1(n57[4]));   // g:/fpga/mxo2/system/project/baud_generator.v(20[10:20])
    defparam cnt_1985_add_4_5.INIT0 = 16'hfaaa;
    defparam cnt_1985_add_4_5.INIT1 = 16'hfaaa;
    defparam cnt_1985_add_4_5.INJECT1_0 = "NO";
    defparam cnt_1985_add_4_5.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_68 (.A(n23123), .B(cnt[6]), .C(cnt[0]), .D(cnt[4]), 
         .Z(n5)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;
    defparam i1_4_lut_adj_68.init = 16'hccc8;
    CCU2D cnt_1985_add_4_3 (.A0(cnt[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n20555), 
          .COUT(n20556), .S0(n57[1]), .S1(n57[2]));   // g:/fpga/mxo2/system/project/baud_generator.v(20[10:20])
    defparam cnt_1985_add_4_3.INIT0 = 16'hfaaa;
    defparam cnt_1985_add_4_3.INIT1 = 16'hfaaa;
    defparam cnt_1985_add_4_3.INJECT1_0 = "NO";
    defparam cnt_1985_add_4_3.INJECT1_1 = "NO";
    LUT4 i2_2_lut (.A(cnt[7]), .B(cnt[5]), .Z(n6)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2_2_lut.init = 16'h8888;
    CCU2D cnt_1985_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n20555), .S1(n57[0]));   // g:/fpga/mxo2/system/project/baud_generator.v(20[10:20])
    defparam cnt_1985_add_4_1.INIT0 = 16'hF000;
    defparam cnt_1985_add_4_1.INIT1 = 16'h0555;
    defparam cnt_1985_add_4_1.INJECT1_0 = "NO";
    defparam cnt_1985_add_4_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module baud_generator_U0
//

module baud_generator_U0 (bps_clk_rx, clk_c, bps_en_rx, GND_net) /* synthesis syn_module_defined=1 */ ;
    output bps_clk_rx;
    input clk_c;
    input bps_en_rx;
    input GND_net;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // g:/fpga/mxo2/system/project/system_top.v(2[15:18])
    
    wire bps_clk_N_2900;
    wire [12:0]cnt;   // g:/fpga/mxo2/system/project/baud_generator.v(12[15:18])
    
    wire cnt_12__N_2896;
    wire [12:0]n57;
    
    wire n7, n23630, n8, n23120, n25736, n20807, n5, n6, n20553, 
        n20552, n20551, n20550, n20549, n20548;
    
    FD1S3AX bps_clk_17 (.D(bps_clk_N_2900), .CK(clk_c), .Q(bps_clk_rx)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=1, LSE_RCOL=2, LSE_LLINE=114, LSE_RLINE=120 */ ;   // g:/fpga/mxo2/system/project/baud_generator.v(28[8] 31[20])
    defparam bps_clk_17.GSR = "ENABLED";
    FD1S3IX cnt_1983__i0 (.D(n57[0]), .CK(clk_c), .CD(cnt_12__N_2896), 
            .Q(cnt[0])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/baud_generator.v(20[10:20])
    defparam cnt_1983__i0.GSR = "ENABLED";
    LUT4 i21460_4_lut (.A(cnt[0]), .B(n7), .C(cnt[6]), .D(n23630), .Z(bps_clk_N_2900)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // g:/fpga/mxo2/system/project/baud_generator.v(28[11:31])
    defparam i21460_4_lut.init = 16'h2000;
    LUT4 i1_4_lut (.A(cnt[9]), .B(cnt[8]), .C(n8), .D(n23120), .Z(n7)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i1_4_lut.init = 16'hfffd;
    LUT4 i20770_2_lut (.A(cnt[5]), .B(cnt[4]), .Z(n23630)) /* synthesis lut_function=(A (B)) */ ;
    defparam i20770_2_lut.init = 16'h8888;
    LUT4 i2_3_lut (.A(cnt[1]), .B(cnt[2]), .C(cnt[3]), .Z(n23120)) /* synthesis lut_function=(A+(B+(C))) */ ;   // g:/fpga/mxo2/system/project/baud_generator.v(17[10:40])
    defparam i2_3_lut.init = 16'hfefe;
    FD1S3IX cnt_1983__i1 (.D(n57[1]), .CK(clk_c), .CD(cnt_12__N_2896), 
            .Q(cnt[1])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/baud_generator.v(20[10:20])
    defparam cnt_1983__i1.GSR = "ENABLED";
    FD1S3IX cnt_1983__i2 (.D(n57[2]), .CK(clk_c), .CD(cnt_12__N_2896), 
            .Q(cnt[2])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/baud_generator.v(20[10:20])
    defparam cnt_1983__i2.GSR = "ENABLED";
    FD1S3IX cnt_1983__i3 (.D(n57[3]), .CK(clk_c), .CD(cnt_12__N_2896), 
            .Q(cnt[3])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/baud_generator.v(20[10:20])
    defparam cnt_1983__i3.GSR = "ENABLED";
    FD1S3IX cnt_1983__i4 (.D(n57[4]), .CK(clk_c), .CD(cnt_12__N_2896), 
            .Q(cnt[4])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/baud_generator.v(20[10:20])
    defparam cnt_1983__i4.GSR = "ENABLED";
    FD1S3IX cnt_1983__i5 (.D(n57[5]), .CK(clk_c), .CD(cnt_12__N_2896), 
            .Q(cnt[5])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/baud_generator.v(20[10:20])
    defparam cnt_1983__i5.GSR = "ENABLED";
    FD1S3IX cnt_1983__i6 (.D(n57[6]), .CK(clk_c), .CD(cnt_12__N_2896), 
            .Q(cnt[6])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/baud_generator.v(20[10:20])
    defparam cnt_1983__i6.GSR = "ENABLED";
    FD1S3IX cnt_1983__i7 (.D(n57[7]), .CK(clk_c), .CD(cnt_12__N_2896), 
            .Q(cnt[7])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/baud_generator.v(20[10:20])
    defparam cnt_1983__i7.GSR = "ENABLED";
    FD1S3IX cnt_1983__i8 (.D(n57[8]), .CK(clk_c), .CD(cnt_12__N_2896), 
            .Q(cnt[8])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/baud_generator.v(20[10:20])
    defparam cnt_1983__i8.GSR = "ENABLED";
    FD1S3IX cnt_1983__i9 (.D(n57[9]), .CK(clk_c), .CD(cnt_12__N_2896), 
            .Q(cnt[9])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/baud_generator.v(20[10:20])
    defparam cnt_1983__i9.GSR = "ENABLED";
    FD1S3IX cnt_1983__i10 (.D(n57[10]), .CK(clk_c), .CD(cnt_12__N_2896), 
            .Q(cnt[10])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/baud_generator.v(20[10:20])
    defparam cnt_1983__i10.GSR = "ENABLED";
    FD1S3IX cnt_1983__i11 (.D(n57[11]), .CK(clk_c), .CD(cnt_12__N_2896), 
            .Q(cnt[11])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/baud_generator.v(20[10:20])
    defparam cnt_1983__i11.GSR = "ENABLED";
    FD1S3IX cnt_1983__i12 (.D(n57[12]), .CK(clk_c), .CD(cnt_12__N_2896), 
            .Q(cnt[12])) /* synthesis syn_use_carry_chain=1 */ ;   // g:/fpga/mxo2/system/project/baud_generator.v(20[10:20])
    defparam cnt_1983__i12.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_454 (.A(cnt[12]), .B(cnt[11]), .Z(n25736)) /* synthesis lut_function=(A+(B)) */ ;   // g:/fpga/mxo2/system/project/baud_generator.v(17[10:40])
    defparam i1_2_lut_rep_454.init = 16'heeee;
    LUT4 i3_3_lut_4_lut (.A(cnt[12]), .B(cnt[11]), .C(cnt[10]), .D(cnt[7]), 
         .Z(n8)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // g:/fpga/mxo2/system/project/baud_generator.v(17[10:40])
    defparam i3_3_lut_4_lut.init = 16'hfffe;
    LUT4 i2_4_lut (.A(n25736), .B(n20807), .C(bps_en_rx), .D(cnt[10]), 
         .Z(cnt_12__N_2896)) /* synthesis lut_function=(A+(B ((D)+!C)+!B !(C))) */ ;   // g:/fpga/mxo2/system/project/baud_generator.v(17[10:40])
    defparam i2_4_lut.init = 16'hefaf;
    LUT4 i2_4_lut_adj_65 (.A(cnt[9]), .B(cnt[8]), .C(n5), .D(n6), .Z(n20807)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_65.init = 16'hfeee;
    LUT4 i1_4_lut_adj_66 (.A(n23120), .B(cnt[6]), .C(cnt[0]), .D(cnt[4]), 
         .Z(n5)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;
    defparam i1_4_lut_adj_66.init = 16'hccc8;
    LUT4 i2_2_lut (.A(cnt[7]), .B(cnt[5]), .Z(n6)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2_2_lut.init = 16'h8888;
    CCU2D cnt_1983_add_4_13 (.A0(cnt[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n20553), .S0(n57[11]), .S1(n57[12]));   // g:/fpga/mxo2/system/project/baud_generator.v(20[10:20])
    defparam cnt_1983_add_4_13.INIT0 = 16'hfaaa;
    defparam cnt_1983_add_4_13.INIT1 = 16'hfaaa;
    defparam cnt_1983_add_4_13.INJECT1_0 = "NO";
    defparam cnt_1983_add_4_13.INJECT1_1 = "NO";
    CCU2D cnt_1983_add_4_11 (.A0(cnt[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n20552), .COUT(n20553), .S0(n57[9]), .S1(n57[10]));   // g:/fpga/mxo2/system/project/baud_generator.v(20[10:20])
    defparam cnt_1983_add_4_11.INIT0 = 16'hfaaa;
    defparam cnt_1983_add_4_11.INIT1 = 16'hfaaa;
    defparam cnt_1983_add_4_11.INJECT1_0 = "NO";
    defparam cnt_1983_add_4_11.INJECT1_1 = "NO";
    CCU2D cnt_1983_add_4_9 (.A0(cnt[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n20551), 
          .COUT(n20552), .S0(n57[7]), .S1(n57[8]));   // g:/fpga/mxo2/system/project/baud_generator.v(20[10:20])
    defparam cnt_1983_add_4_9.INIT0 = 16'hfaaa;
    defparam cnt_1983_add_4_9.INIT1 = 16'hfaaa;
    defparam cnt_1983_add_4_9.INJECT1_0 = "NO";
    defparam cnt_1983_add_4_9.INJECT1_1 = "NO";
    CCU2D cnt_1983_add_4_7 (.A0(cnt[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n20550), 
          .COUT(n20551), .S0(n57[5]), .S1(n57[6]));   // g:/fpga/mxo2/system/project/baud_generator.v(20[10:20])
    defparam cnt_1983_add_4_7.INIT0 = 16'hfaaa;
    defparam cnt_1983_add_4_7.INIT1 = 16'hfaaa;
    defparam cnt_1983_add_4_7.INJECT1_0 = "NO";
    defparam cnt_1983_add_4_7.INJECT1_1 = "NO";
    CCU2D cnt_1983_add_4_5 (.A0(cnt[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n20549), 
          .COUT(n20550), .S0(n57[3]), .S1(n57[4]));   // g:/fpga/mxo2/system/project/baud_generator.v(20[10:20])
    defparam cnt_1983_add_4_5.INIT0 = 16'hfaaa;
    defparam cnt_1983_add_4_5.INIT1 = 16'hfaaa;
    defparam cnt_1983_add_4_5.INJECT1_0 = "NO";
    defparam cnt_1983_add_4_5.INJECT1_1 = "NO";
    CCU2D cnt_1983_add_4_3 (.A0(cnt[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n20548), 
          .COUT(n20549), .S0(n57[1]), .S1(n57[2]));   // g:/fpga/mxo2/system/project/baud_generator.v(20[10:20])
    defparam cnt_1983_add_4_3.INIT0 = 16'hfaaa;
    defparam cnt_1983_add_4_3.INIT1 = 16'hfaaa;
    defparam cnt_1983_add_4_3.INJECT1_0 = "NO";
    defparam cnt_1983_add_4_3.INJECT1_1 = "NO";
    CCU2D cnt_1983_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n20548), .S1(n57[0]));   // g:/fpga/mxo2/system/project/baud_generator.v(20[10:20])
    defparam cnt_1983_add_4_1.INIT0 = 16'hF000;
    defparam cnt_1983_add_4_1.INIT1 = 16'h0555;
    defparam cnt_1983_add_4_1.INJECT1_0 = "NO";
    defparam cnt_1983_add_4_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module DS18B20Z
//

module DS18B20Z (clk_1mhz, clk_c, \tamp_data[0] , clk_c_enable_931, 
            tamp_out_11__N_495, \state_back_2__N_261[2] , one_wire_N_501, 
            \state[0] , clk_c_enable_1439, \data_out[0] , \cnt_read[2] , 
            \state[1] , \tamp_data[9] , \tamp_data[8] , \tamp_data[7] , 
            \tamp_data[6] , \tamp_data[5] , \tamp_data[4] , \tamp_data[2] , 
            tamp_out_11__N_483, \tamp_data[1] , tamp_out_11__N_489, clk_c_enable_686, 
            clk_c_enable_117, clk_c_enable_132, one_wire_out, n25765, 
            n50, GND_net, n25618, n25607, clk_c_enable_684, \num_delay_19__N_369[5] , 
            clk_c_enable_688, \data_out[1] , \data_out[2] , \tamp_out_11__N_478[3] , 
            \tamp_data[3] , n20945, \cnt_init[2] , n25689, clk_c_enable_1433, 
            clk_c_enable_1437, n23656, n28, n16451, n16602, n25742, 
            n5709, n37, n29, n25484, n25453, n25857) /* synthesis syn_module_defined=1 */ ;
    output clk_1mhz;
    input clk_c;
    output \tamp_data[0] ;
    input clk_c_enable_931;
    input tamp_out_11__N_495;
    output \state_back_2__N_261[2] ;
    output one_wire_N_501;
    output \state[0] ;
    input clk_c_enable_1439;
    output \data_out[0] ;
    output \cnt_read[2] ;
    output \state[1] ;
    output \tamp_data[9] ;
    output \tamp_data[8] ;
    output \tamp_data[7] ;
    output \tamp_data[6] ;
    output \tamp_data[5] ;
    output \tamp_data[4] ;
    output \tamp_data[2] ;
    input tamp_out_11__N_483;
    output \tamp_data[1] ;
    input tamp_out_11__N_489;
    input clk_c_enable_686;
    input clk_c_enable_117;
    input clk_c_enable_132;
    input one_wire_out;
    output n25765;
    output n50;
    input GND_net;
    input n25618;
    input n25607;
    input clk_c_enable_684;
    input \num_delay_19__N_369[5] ;
    input clk_c_enable_688;
    output \data_out[1] ;
    output \data_out[2] ;
    output \tamp_out_11__N_478[3] ;
    output \tamp_data[3] ;
    input n20945;
    output \cnt_init[2] ;
    output n25689;
    input clk_c_enable_1433;
    input clk_c_enable_1437;
    input n23656;
    output n28;
    output n16451;
    output n16602;
    output n25742;
    output n5709;
    output n37;
    output n29;
    output n25484;
    output n25453;
    output n25857;
    
    wire clk_1mhz /* synthesis is_clock=1, SET_AS_NETWORK=\DS18B20Z_inst/clk_1mhz */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(18[9:17])
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // g:/fpga/mxo2/system/project/system_top.v(2[15:18])
    
    wire clk_1mhz_N_503;
    wire [3:0]cnt_write;   // g:/fpga/mxo2/system/project/ds18b20z.v(40[13:22])
    
    wire n5035;
    wire [3:0]cnt_write_3__N_333;
    
    wire n329;
    wire [19:0]n331;
    wire [19:0]cnt_delay_19__N_187;
    
    wire one_wire_N_504, n2, n3, n23827, one_wire_N_515, n13, n14, 
        one_wire_N_510;
    wire [2:0]cnt_read;   // g:/fpga/mxo2/system/project/ds18b20z.v(41[13:21])
    wire [2:0]state_back;   // g:/fpga/mxo2/system/project/ds18b20z.v(45[14:24])
    
    wire n4, n7;
    wire [2:0]cnt;   // g:/fpga/mxo2/system/project/ds18b20z.v(32[13:16])
    wire [2:0]cnt_2__N_161;
    
    wire n25680, n25627, n32, clk_c_enable_748;
    wire [15:0]temperature;   // g:/fpga/mxo2/system/project/ds18b20z.v(42[14:25])
    
    wire clk_c_enable_709;
    wire [7:0]temperature_buffer;   // g:/fpga/mxo2/system/project/ds18b20z.v(43[13:31])
    
    wire clk_c_enable_717;
    wire [19:0]cnt_delay;   // g:/fpga/mxo2/system/project/ds18b20z.v(38[14:23])
    
    wire clk_c_enable_736, n23294, clk_c_enable_26;
    wire [2:0]state_back_2__N_261;
    
    wire n23814, n25448, n25850, n25851;
    wire [6:0]n1854;
    wire [8:0]data_out;   // g:/fpga/mxo2/system/project/ds18b20z.v(46[20:28])
    wire [7:0]data_wr;   // g:/fpga/mxo2/system/project/ds18b20z.v(35[13:20])
    
    wire clk_c_enable_83, n7_adj_5022, n7_adj_5023, n25717;
    wire [7:0]data_wr_buffer;   // g:/fpga/mxo2/system/project/ds18b20z.v(36[13:27])
    
    wire clk_c_enable_86, n25452;
    wire [19:0]num_delay;   // g:/fpga/mxo2/system/project/ds18b20z.v(39[14:23])
    wire [19:0]num_delay_19__N_369;
    wire [2:0]state_2__N_258;
    
    wire clk_c_enable_201;
    wire [3:0]cnt_main;   // g:/fpga/mxo2/system/project/ds18b20z.v(34[13:21])
    
    wire n25477, n25476, clk_c_enable_614, n25687;
    wire [2:0]state_2__N_306;
    wire [2:0]state_2__N_303;
    
    wire n2_adj_5024, n16018, n4_adj_5025, clk_c_enable_545, clk_c_enable_553, 
        clk_c_enable_557, n14912, n21141, n14920, n25775, n25776, 
        clk_c_enable_1416, clk_c_enable_634;
    wire [2:0]cnt_1mhz;   // g:/fpga/mxo2/system/project/ds18b20z.v(19[13:21])
    wire [2:0]n17;
    
    wire n25741, n25584, n20481, n20482, n25626, n25705, n25449, 
        n25669, n25478, n25480, n25739, n12075, n15869, one_wire_N_502, 
        n25852, n25853, clk_c_enable_683, clk_c_enable_1420, n12080, 
        n25668, n25722, n44, n23162, n23481, clk_c_enable_1372, 
        n20667, clk_c_enable_689, n25740, n25475, n25708, n23114;
    wire [3:0]tamp_out_11__N_414;
    
    wire n25013, n25591, n25592, clk_c_enable_747, n25679, n30, 
        n24034, clk_c_enable_1426, n15328, n25652, n25655, n24678;
    wire [2:0]cnt_init;   // g:/fpga/mxo2/system/project/ds18b20z.v(37[13:21])
    
    wire n1, n2_adj_5026;
    wire [2:0]n253;
    
    wire n23255, clk_c_enable_1422, n25707, n25855, n26776, n25757, 
        n25625, n20480, n20479, n25766, n25767, n24679, n25699, 
        n20584, clk_c_enable_1447;
    wire [2:0]n102;
    
    wire n20583, n20582;
    wire [2:0]n1853;
    
    wire clk_c_enable_1371, n20581, n20580, n20579, n9, n20578, 
        n20577, n20576, n20575, n20_adj_5027, one_wire_N_508, one_wire_N_505, 
        n25663, n25723, n25670, n23372, n23154, n25688, n25644, 
        n3_adj_5028, n2_adj_5029, n8250, n24052, n25450;
    wire [3:0]n25;
    
    wire n6, n14905, n25700, n49, n33, n23436, n3_adj_5030, n21171, 
        n15797, n34, n25451, n23622, n46, n25738, n20488, n25613, 
        n20483, n20484, n25482, n66, n25483, n20487, n20485, n20486, 
        n24036;
    
    FD1S3AX clk_1mhz_194 (.D(clk_1mhz_N_503), .CK(clk_c), .Q(clk_1mhz)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(24[14] 29[8])
    defparam clk_1mhz_194.GSR = "ENABLED";
    LUT4 i20662_3_lut_4_lut (.A(cnt_write[0]), .B(cnt_write[1]), .C(cnt_write[2]), 
         .D(n5035), .Z(cnt_write_3__N_333[2])) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(115[30] 118[24])
    defparam i20662_3_lut_4_lut.init = 16'h0078;
    FD1P3AX tamp_out__i1 (.D(tamp_out_11__N_495), .SP(clk_c_enable_931), 
            .CK(clk_c), .Q(\tamp_data[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(173[10] 202[8])
    defparam tamp_out__i1.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut (.A(\state_back_2__N_261[2] ), .B(n329), .C(n331[12]), 
         .Z(cnt_delay_19__N_187[12])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut.init = 16'h2020;
    FD1S3AX one_wire_buffer_204 (.D(one_wire_N_504), .CK(clk_1mhz), .Q(one_wire_N_501)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam one_wire_buffer_204.GSR = "ENABLED";
    PFUMX state_2__I_0_i7 (.BLUT(n2), .ALUT(n3), .C0(n23827), .Z(one_wire_N_515)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;
    PFUMX i16 (.BLUT(n13), .ALUT(n14), .C0(n23827), .Z(one_wire_N_510));
    LUT4 i11_4_lut (.A(cnt_read[1]), .B(state_back[0]), .C(\state[0] ), 
         .D(n4), .Z(n7)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B+!(C))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(44[14:19])
    defparam i11_4_lut.init = 16'hc5cf;
    FD1P3AX cnt_i0_i0 (.D(cnt_2__N_161[0]), .SP(clk_c_enable_1439), .CK(clk_c), 
            .Q(cnt[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam cnt_i0_i0.GSR = "ENABLED";
    LUT4 i1_3_lut_4_lut (.A(n25680), .B(n25627), .C(n32), .D(\state_back_2__N_261[2] ), 
         .Z(clk_c_enable_748)) /* synthesis lut_function=(!(A+!(B (C+(D))))) */ ;
    defparam i1_3_lut_4_lut.init = 16'h4440;
    FD1P3AX temperature_i0_i0 (.D(temperature_buffer[0]), .SP(clk_c_enable_709), 
            .CK(clk_c), .Q(temperature[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam temperature_i0_i0.GSR = "ENABLED";
    FD1P3AX data_out_i0_i0 (.D(temperature[0]), .SP(clk_c_enable_717), .CK(clk_c), 
            .Q(\data_out[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam data_out_i0_i0.GSR = "ENABLED";
    FD1P3AX cnt_delay_i0_i0 (.D(n23294), .SP(clk_c_enable_736), .CK(clk_c), 
            .Q(cnt_delay[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam cnt_delay_i0_i0.GSR = "ENABLED";
    FD1P3AX state_back_i0_i0 (.D(state_back_2__N_261[0]), .SP(clk_c_enable_26), 
            .CK(clk_c), .Q(state_back[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam state_back_i0_i0.GSR = "ENABLED";
    LUT4 n23814_bdd_4_lut (.A(n23814), .B(\cnt_read[2] ), .C(\state[0] ), 
         .D(\state[1] ), .Z(n25448)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam n23814_bdd_4_lut.init = 16'hfff7;
    LUT4 n25850_bdd_2_lut (.A(n25850), .B(\state_back_2__N_261[2] ), .Z(n25851)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam n25850_bdd_2_lut.init = 16'h2222;
    FD1P3AX tamp_out__i10 (.D(n1854[5]), .SP(clk_c_enable_931), .CK(clk_c), 
            .Q(\tamp_data[9] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(173[10] 202[8])
    defparam tamp_out__i10.GSR = "ENABLED";
    FD1P3AX tamp_out__i9 (.D(n1854[4]), .SP(clk_c_enable_931), .CK(clk_c), 
            .Q(\tamp_data[8] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(173[10] 202[8])
    defparam tamp_out__i9.GSR = "ENABLED";
    FD1P3AX tamp_out__i8 (.D(n1854[3]), .SP(clk_c_enable_931), .CK(clk_c), 
            .Q(\tamp_data[7] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(173[10] 202[8])
    defparam tamp_out__i8.GSR = "ENABLED";
    FD1P3AX tamp_out__i7 (.D(n1854[2]), .SP(clk_c_enable_931), .CK(clk_c), 
            .Q(\tamp_data[6] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(173[10] 202[8])
    defparam tamp_out__i7.GSR = "ENABLED";
    FD1P3AX tamp_out__i6 (.D(n1854[1]), .SP(clk_c_enable_931), .CK(clk_c), 
            .Q(\tamp_data[5] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(173[10] 202[8])
    defparam tamp_out__i6.GSR = "ENABLED";
    FD1P3AX tamp_out__i5 (.D(data_out[4]), .SP(clk_c_enable_931), .CK(clk_c), 
            .Q(\tamp_data[4] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(173[10] 202[8])
    defparam tamp_out__i5.GSR = "ENABLED";
    FD1P3AX tamp_out__i3 (.D(tamp_out_11__N_483), .SP(clk_c_enable_931), 
            .CK(clk_c), .Q(\tamp_data[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(173[10] 202[8])
    defparam tamp_out__i3.GSR = "ENABLED";
    FD1P3AX tamp_out__i2 (.D(tamp_out_11__N_489), .SP(clk_c_enable_931), 
            .CK(clk_c), .Q(\tamp_data[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(173[10] 202[8])
    defparam tamp_out__i2.GSR = "ENABLED";
    FD1P3AX data_wr_i0_i7 (.D(n7_adj_5022), .SP(clk_c_enable_83), .CK(clk_c), 
            .Q(data_wr[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam data_wr_i0_i7.GSR = "DISABLED";
    FD1P3AX data_wr_i0_i6 (.D(n7_adj_5023), .SP(clk_c_enable_83), .CK(clk_c), 
            .Q(data_wr[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam data_wr_i0_i6.GSR = "DISABLED";
    FD1P3AX data_wr_i0_i1 (.D(n25717), .SP(clk_c_enable_83), .CK(clk_c), 
            .Q(data_wr[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam data_wr_i0_i1.GSR = "DISABLED";
    FD1P3AX data_wr_buffer_i0_i7 (.D(data_wr[7]), .SP(clk_c_enable_86), 
            .CK(clk_c), .Q(data_wr_buffer[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam data_wr_buffer_i0_i7.GSR = "DISABLED";
    FD1P3AX data_wr_buffer_i0_i6 (.D(data_wr[6]), .SP(clk_c_enable_86), 
            .CK(clk_c), .Q(data_wr_buffer[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam data_wr_buffer_i0_i6.GSR = "DISABLED";
    FD1P3AX data_wr_buffer_i0_i4 (.D(data_wr[1]), .SP(clk_c_enable_86), 
            .CK(clk_c), .Q(data_wr_buffer[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam data_wr_buffer_i0_i4.GSR = "DISABLED";
    LUT4 n5035_bdd_3_lut_22454 (.A(n5035), .B(\state[0] ), .C(\state[1] ), 
         .Z(n25452)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B+(C))) */ ;
    defparam n5035_bdd_3_lut_22454.init = 16'h8383;
    FD1P3AX num_delay_i0_i0 (.D(num_delay_19__N_369[0]), .SP(clk_c_enable_686), 
            .CK(clk_c), .Q(num_delay[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam num_delay_i0_i0.GSR = "DISABLED";
    FD1P3AX num_delay_i0_i2 (.D(num_delay_19__N_369[2]), .SP(clk_c_enable_117), 
            .CK(clk_c), .Q(num_delay[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam num_delay_i0_i2.GSR = "DISABLED";
    FD1P3AX state_i0_i0 (.D(state_2__N_258[0]), .SP(clk_c_enable_132), .CK(clk_c), 
            .Q(\state[0] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam state_i0_i0.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_adj_19 (.A(\state_back_2__N_261[2] ), .B(n329), 
         .C(n331[13]), .Z(cnt_delay_19__N_187[13])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_19.init = 16'h2020;
    FD1P3AX temperature_buffer_i0_i1 (.D(one_wire_out), .SP(clk_c_enable_201), 
            .CK(clk_c), .Q(temperature_buffer[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam temperature_buffer_i0_i1.GSR = "DISABLED";
    LUT4 cnt_main_2__bdd_4_lut (.A(cnt_main[2]), .B(cnt_main[1]), .C(cnt_main[3]), 
         .D(cnt_main[0]), .Z(n25477)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (B (C+!(D))+!B !(C (D))))) */ ;
    defparam cnt_main_2__bdd_4_lut.init = 16'h1c00;
    LUT4 cnt_main_2__bdd_1_lut (.A(cnt_write[3]), .Z(n25476)) /* synthesis lut_function=(!(A)) */ ;
    defparam cnt_main_2__bdd_1_lut.init = 16'h5555;
    FD1P3AX num_delay_i0_i12 (.D(n25687), .SP(clk_c_enable_614), .CK(clk_c), 
            .Q(num_delay[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam num_delay_i0_i12.GSR = "DISABLED";
    LUT4 i1_2_lut_3_lut_adj_20 (.A(\state_back_2__N_261[2] ), .B(n329), 
         .C(n331[14]), .Z(cnt_delay_19__N_187[14])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_20.init = 16'h2020;
    PFUMX state_2__I_0_216_Mux_0_i2 (.BLUT(state_2__N_306[0]), .ALUT(state_2__N_303[0]), 
          .C0(\state[0] ), .Z(n2_adj_5024)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;
    LUT4 state_2__I_0_i3_4_lut (.A(\state[0] ), .B(n16018), .C(\state_back_2__N_261[2] ), 
         .D(n4_adj_5025), .Z(n3)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(62[9] 163[16])
    defparam state_2__I_0_i3_4_lut.init = 16'hfaca;
    LUT4 i1_2_lut_3_lut_adj_21 (.A(\state_back_2__N_261[2] ), .B(n329), 
         .C(n331[15]), .Z(cnt_delay_19__N_187[15])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_21.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_22 (.A(\state_back_2__N_261[2] ), .B(n329), 
         .C(n331[6]), .Z(cnt_delay_19__N_187[6])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_22.init = 16'h2020;
    FD1P3AX temperature_buffer_i0_i2 (.D(one_wire_out), .SP(clk_c_enable_545), 
            .CK(clk_c), .Q(temperature_buffer[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam temperature_buffer_i0_i2.GSR = "DISABLED";
    FD1P3AX temperature_buffer_i0_i3 (.D(one_wire_out), .SP(clk_c_enable_553), 
            .CK(clk_c), .Q(temperature_buffer[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam temperature_buffer_i0_i3.GSR = "DISABLED";
    FD1P3AX temperature_buffer_i0_i4 (.D(one_wire_out), .SP(clk_c_enable_557), 
            .CK(clk_c), .Q(temperature_buffer[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam temperature_buffer_i0_i4.GSR = "DISABLED";
    PFUMX i12127 (.BLUT(n14912), .ALUT(n21141), .C0(\state[1] ), .Z(n14920));
    PFUMX i22157 (.BLUT(n25775), .ALUT(n25776), .C0(\state[1] ), .Z(clk_c_enable_1416));
    FD1P3AX num_delay_i0_i8 (.D(num_delay_19__N_369[8]), .SP(clk_c_enable_614), 
            .CK(clk_c), .Q(num_delay[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam num_delay_i0_i8.GSR = "DISABLED";
    FD1P3AX temperature_buffer_i0_i5 (.D(one_wire_out), .SP(clk_c_enable_634), 
            .CK(clk_c), .Q(temperature_buffer[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam temperature_buffer_i0_i5.GSR = "DISABLED";
    FD1S3IX cnt_1mhz_1980__i0 (.D(n17[0]), .CK(clk_c), .CD(n25765), .Q(cnt_1mhz[0]));   // g:/fpga/mxo2/system/project/ds18b20z.v(28[21:36])
    defparam cnt_1mhz_1980__i0.GSR = "ENABLED";
    LUT4 i1_3_lut_4_lut_4_lut (.A(n25741), .B(n25627), .C(n50), .D(n25584), 
         .Z(clk_c_enable_614)) /* synthesis lut_function=(A (B (C (D)))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(44[14:19])
    defparam i1_3_lut_4_lut_4_lut.init = 16'hc040;
    CCU2D add_76_7 (.A0(cnt_delay[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt_delay[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n20481), .COUT(n20482), .S0(n331[5]), .S1(n331[6]));   // g:/fpga/mxo2/system/project/ds18b20z.v(161[43:59])
    defparam add_76_7.INIT0 = 16'h5aaa;
    defparam add_76_7.INIT1 = 16'h5aaa;
    defparam add_76_7.INJECT1_0 = "NO";
    defparam add_76_7.INJECT1_1 = "NO";
    LUT4 i1_3_lut_4_lut_4_lut_adj_23 (.A(n25687), .B(n25618), .C(n25626), 
         .D(\state[0] ), .Z(n50)) /* synthesis lut_function=(A (B (C (D)))+!A (B)) */ ;
    defparam i1_3_lut_4_lut_4_lut_adj_23.init = 16'hc444;
    LUT4 n23814_bdd_3_lut_4_lut (.A(n25705), .B(cnt_write[3]), .C(\state[1] ), 
         .D(\state[0] ), .Z(n25449)) /* synthesis lut_function=(!(A (C (D))+!A (B (C (D))))) */ ;
    defparam n23814_bdd_3_lut_4_lut.init = 16'h1fff;
    LUT4 n25479_bdd_3_lut_4_lut (.A(n25669), .B(\state[1] ), .C(\state[0] ), 
         .D(n25478), .Z(n25480)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;
    defparam n25479_bdd_3_lut_4_lut.init = 16'hf808;
    LUT4 i9260_3_lut_4_lut (.A(\state[0] ), .B(n25607), .C(\state[1] ), 
         .D(n25739), .Z(n12075)) /* synthesis lut_function=(!(A+(B+!((D)+!C)))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam i9260_3_lut_4_lut.init = 16'h1101;
    LUT4 i21346_2_lut_4_lut (.A(\cnt_read[2] ), .B(\state_back_2__N_261[2] ), 
         .C(n23814), .D(cnt_read[0]), .Z(n15869)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A ((D)+!B))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(62[9] 163[16])
    defparam i21346_2_lut_4_lut.init = 16'h004c;
    FD1P3AX i136_211 (.D(one_wire_N_515), .SP(one_wire_N_510), .CK(clk_1mhz), 
            .Q(one_wire_N_502)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam i136_211.GSR = "ENABLED";
    PFUMX i22204 (.BLUT(n25852), .ALUT(n25851), .C0(\state[1] ), .Z(n25853));
    FD1P3AX num_delay_i0_i6 (.D(num_delay_19__N_369[6]), .SP(clk_c_enable_683), 
            .CK(clk_c), .Q(num_delay[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam num_delay_i0_i6.GSR = "DISABLED";
    LUT4 i9265_2_lut_4_lut (.A(\cnt_read[2] ), .B(\state_back_2__N_261[2] ), 
         .C(n23814), .D(clk_c_enable_1420), .Z(n12080)) /* synthesis lut_function=(A (B (C (D))+!B (D))+!A !(B+!(D))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(62[9] 163[16])
    defparam i9265_2_lut_4_lut.init = 16'hb300;
    FD1P3AX num_delay_i0_i5 (.D(\num_delay_19__N_369[5] ), .SP(clk_c_enable_684), 
            .CK(clk_c), .Q(num_delay[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam num_delay_i0_i5.GSR = "DISABLED";
    LUT4 i1_4_lut (.A(cnt_write[3]), .B(\state_back_2__N_261[2] ), .C(n25668), 
         .D(n25722), .Z(n44)) /* synthesis lut_function=(A (B)+!A (B+(C (D)))) */ ;
    defparam i1_4_lut.init = 16'hdccc;
    LUT4 i21538_4_lut (.A(n25680), .B(n23162), .C(\state_back_2__N_261[2] ), 
         .D(n23481), .Z(clk_c_enable_1372)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;
    defparam i21538_4_lut.init = 16'h1011;
    LUT4 i17_4_lut (.A(n14920), .B(n20667), .C(\state_back_2__N_261[2] ), 
         .D(\state[1] ), .Z(state_2__N_258[1])) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(44[14:19])
    defparam i17_4_lut.init = 16'hfaca;
    LUT4 i1_2_lut_4_lut (.A(n25722), .B(cnt_write[3]), .C(\state_back_2__N_261[2] ), 
         .D(n25668), .Z(n23162)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(62[9] 163[16])
    defparam i1_2_lut_4_lut.init = 16'h0200;
    LUT4 i2_3_lut (.A(state_back[1]), .B(\state[0] ), .C(n329), .Z(n20667)) /* synthesis lut_function=(A (B (C))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(44[14:19])
    defparam i2_3_lut.init = 16'h8080;
    FD1P3AX num_delay_i0_i4 (.D(num_delay_19__N_369[4]), .SP(clk_c_enable_688), 
            .CK(clk_c), .Q(num_delay[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam num_delay_i0_i4.GSR = "DISABLED";
    FD1P3AX num_delay_i0_i3 (.D(num_delay_19__N_369[3]), .SP(clk_c_enable_686), 
            .CK(clk_c), .Q(num_delay[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam num_delay_i0_i3.GSR = "DISABLED";
    FD1P3AX num_delay_i0_i1 (.D(num_delay_19__N_369[1]), .SP(clk_c_enable_688), 
            .CK(clk_c), .Q(num_delay[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam num_delay_i0_i1.GSR = "DISABLED";
    FD1P3AX temperature_buffer_i0_i6 (.D(one_wire_out), .SP(clk_c_enable_689), 
            .CK(clk_c), .Q(temperature_buffer[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam temperature_buffer_i0_i6.GSR = "DISABLED";
    LUT4 n8345_bdd_3_lut_4_lut (.A(cnt_read[0]), .B(n25740), .C(state_back[2]), 
         .D(\state[0] ), .Z(n25475)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C (D))) */ ;
    defparam n8345_bdd_3_lut_4_lut.init = 16'hf022;
    LUT4 i1_3_lut_rep_345_4_lut (.A(cnt_read[0]), .B(n25740), .C(\state_back_2__N_261[2] ), 
         .D(n25708), .Z(n25627)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (C))) */ ;
    defparam i1_3_lut_rep_345_4_lut.init = 16'h0f2f;
    LUT4 i21365_2_lut_3_lut_4_lut (.A(cnt[1]), .B(n23114), .C(cnt[2]), 
         .D(cnt[0]), .Z(clk_c_enable_545)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i21365_2_lut_3_lut_4_lut.init = 16'h0002;
    FD1P3AX temperature_i0_i1 (.D(temperature_buffer[1]), .SP(clk_c_enable_709), 
            .CK(clk_c), .Q(temperature[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam temperature_i0_i1.GSR = "ENABLED";
    FD1P3AX temperature_i0_i2 (.D(temperature_buffer[2]), .SP(clk_c_enable_709), 
            .CK(clk_c), .Q(temperature[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam temperature_i0_i2.GSR = "ENABLED";
    FD1P3AX temperature_i0_i3 (.D(temperature_buffer[3]), .SP(clk_c_enable_709), 
            .CK(clk_c), .Q(temperature[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam temperature_i0_i3.GSR = "ENABLED";
    FD1P3AX temperature_i0_i4 (.D(temperature_buffer[4]), .SP(clk_c_enable_709), 
            .CK(clk_c), .Q(temperature[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam temperature_i0_i4.GSR = "ENABLED";
    FD1P3AX temperature_i0_i5 (.D(temperature_buffer[5]), .SP(clk_c_enable_709), 
            .CK(clk_c), .Q(temperature[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam temperature_i0_i5.GSR = "ENABLED";
    FD1P3AX temperature_i0_i6 (.D(temperature_buffer[6]), .SP(clk_c_enable_709), 
            .CK(clk_c), .Q(temperature[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam temperature_i0_i6.GSR = "ENABLED";
    FD1P3AX temperature_i0_i7 (.D(temperature_buffer[7]), .SP(clk_c_enable_709), 
            .CK(clk_c), .Q(temperature[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam temperature_i0_i7.GSR = "ENABLED";
    FD1P3AX data_out_i0_i1 (.D(temperature[1]), .SP(clk_c_enable_717), .CK(clk_c), 
            .Q(\data_out[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam data_out_i0_i1.GSR = "ENABLED";
    FD1P3AX data_out_i0_i2 (.D(temperature[2]), .SP(clk_c_enable_717), .CK(clk_c), 
            .Q(\data_out[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam data_out_i0_i2.GSR = "ENABLED";
    FD1P3AX data_out_i0_i3 (.D(temperature[3]), .SP(clk_c_enable_717), .CK(clk_c), 
            .Q(\tamp_out_11__N_478[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam data_out_i0_i3.GSR = "ENABLED";
    FD1P3AX data_out_i0_i4 (.D(temperature[4]), .SP(clk_c_enable_717), .CK(clk_c), 
            .Q(data_out[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam data_out_i0_i4.GSR = "ENABLED";
    FD1P3AX data_out_i0_i5 (.D(temperature[5]), .SP(clk_c_enable_717), .CK(clk_c), 
            .Q(data_out[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam data_out_i0_i5.GSR = "ENABLED";
    FD1P3AX data_out_i0_i6 (.D(temperature[6]), .SP(clk_c_enable_717), .CK(clk_c), 
            .Q(data_out[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam data_out_i0_i6.GSR = "ENABLED";
    FD1P3AX data_out_i0_i7 (.D(temperature[7]), .SP(clk_c_enable_717), .CK(clk_c), 
            .Q(data_out[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam data_out_i0_i7.GSR = "ENABLED";
    FD1P3AX data_out_i0_i8 (.D(temperature[8]), .SP(clk_c_enable_717), .CK(clk_c), 
            .Q(tamp_out_11__N_414[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam data_out_i0_i8.GSR = "ENABLED";
    FD1P3AX cnt_delay_i0_i1 (.D(cnt_delay_19__N_187[1]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(cnt_delay[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam cnt_delay_i0_i1.GSR = "ENABLED";
    FD1P3AX cnt_delay_i0_i2 (.D(cnt_delay_19__N_187[2]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(cnt_delay[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam cnt_delay_i0_i2.GSR = "ENABLED";
    FD1P3AX cnt_delay_i0_i3 (.D(cnt_delay_19__N_187[3]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(cnt_delay[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam cnt_delay_i0_i3.GSR = "ENABLED";
    FD1P3AX cnt_delay_i0_i4 (.D(cnt_delay_19__N_187[4]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(cnt_delay[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam cnt_delay_i0_i4.GSR = "ENABLED";
    FD1P3AX cnt_delay_i0_i5 (.D(cnt_delay_19__N_187[5]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(cnt_delay[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam cnt_delay_i0_i5.GSR = "ENABLED";
    FD1P3AX cnt_delay_i0_i6 (.D(cnt_delay_19__N_187[6]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(cnt_delay[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam cnt_delay_i0_i6.GSR = "ENABLED";
    FD1P3AX cnt_delay_i0_i7 (.D(cnt_delay_19__N_187[7]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(cnt_delay[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam cnt_delay_i0_i7.GSR = "ENABLED";
    FD1P3AX cnt_delay_i0_i8 (.D(cnt_delay_19__N_187[8]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(cnt_delay[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam cnt_delay_i0_i8.GSR = "ENABLED";
    FD1P3AX cnt_delay_i0_i9 (.D(cnt_delay_19__N_187[9]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(cnt_delay[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam cnt_delay_i0_i9.GSR = "ENABLED";
    FD1P3AX cnt_delay_i0_i10 (.D(cnt_delay_19__N_187[10]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(cnt_delay[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam cnt_delay_i0_i10.GSR = "ENABLED";
    FD1P3AX cnt_delay_i0_i11 (.D(cnt_delay_19__N_187[11]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(cnt_delay[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam cnt_delay_i0_i11.GSR = "ENABLED";
    FD1P3AX cnt_delay_i0_i12 (.D(cnt_delay_19__N_187[12]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(cnt_delay[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam cnt_delay_i0_i12.GSR = "ENABLED";
    FD1P3AX cnt_delay_i0_i13 (.D(cnt_delay_19__N_187[13]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(cnt_delay[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam cnt_delay_i0_i13.GSR = "ENABLED";
    FD1P3AX cnt_delay_i0_i14 (.D(cnt_delay_19__N_187[14]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(cnt_delay[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam cnt_delay_i0_i14.GSR = "ENABLED";
    FD1P3AX cnt_delay_i0_i15 (.D(cnt_delay_19__N_187[15]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(cnt_delay[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam cnt_delay_i0_i15.GSR = "ENABLED";
    FD1P3AX cnt_delay_i0_i16 (.D(cnt_delay_19__N_187[16]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(cnt_delay[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam cnt_delay_i0_i16.GSR = "ENABLED";
    FD1P3AX cnt_delay_i0_i17 (.D(cnt_delay_19__N_187[17]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(cnt_delay[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam cnt_delay_i0_i17.GSR = "ENABLED";
    FD1P3AX cnt_delay_i0_i18 (.D(cnt_delay_19__N_187[18]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(cnt_delay[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam cnt_delay_i0_i18.GSR = "ENABLED";
    FD1P3AX cnt_delay_i0_i19 (.D(cnt_delay_19__N_187[19]), .SP(clk_c_enable_736), 
            .CK(clk_c), .Q(cnt_delay[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam cnt_delay_i0_i19.GSR = "ENABLED";
    LUT4 n1058_bdd_2_lut_21821_4_lut_4_lut (.A(n25687), .B(n25013), .C(n25591), 
         .D(n25592), .Z(clk_c_enable_26)) /* synthesis lut_function=(A (B (C (D)))+!A (B (C))) */ ;
    defparam n1058_bdd_2_lut_21821_4_lut_4_lut.init = 16'hc040;
    FD1P3AX temperature_buffer_i0_i7 (.D(one_wire_out), .SP(clk_c_enable_747), 
            .CK(clk_c), .Q(temperature_buffer[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam temperature_buffer_i0_i7.GSR = "DISABLED";
    FD1P3AX state_back_i0_i2 (.D(\state_back_2__N_261[2] ), .SP(clk_c_enable_748), 
            .CK(clk_c), .Q(state_back[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam state_back_i0_i2.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_adj_24 (.A(\state_back_2__N_261[2] ), .B(n329), 
         .C(n331[16]), .Z(cnt_delay_19__N_187[16])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_24.init = 16'h2020;
    LUT4 i1_3_lut_4_lut_adj_25 (.A(cnt_read[0]), .B(n25740), .C(\state_back_2__N_261[2] ), 
         .D(n25679), .Z(n30)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C+(D)))) */ ;
    defparam i1_3_lut_4_lut_adj_25.init = 16'hff10;
    LUT4 i1_4_lut_adj_26 (.A(n25765), .B(clk_1mhz), .C(n24034), .D(\state_back_2__N_261[2] ), 
         .Z(clk_c_enable_1426)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_4_lut_adj_26.init = 16'h0002;
    LUT4 i21319_2_lut (.A(\state[1] ), .B(\state[0] ), .Z(n24034)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i21319_2_lut.init = 16'h6666;
    LUT4 i1_2_lut (.A(\state[1] ), .B(clk_c_enable_1426), .Z(n15328)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut.init = 16'h4444;
    LUT4 i7275_4_lut (.A(cnt_write[0]), .B(n25652), .C(n5035), .D(n25655), 
         .Z(cnt_write_3__N_333[0])) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C)+!B !((D)+!C)))) */ ;
    defparam i7275_4_lut.init = 16'h3505;
    FD1P3IX tamp_out__i4 (.D(\tamp_out_11__N_478[3] ), .SP(clk_c_enable_931), 
            .CD(n20945), .CK(clk_c), .Q(\tamp_data[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(173[10] 202[8])
    defparam tamp_out__i4.GSR = "ENABLED";
    LUT4 i17577_2_lut (.A(cnt_1mhz[1]), .B(cnt_1mhz[0]), .Z(n17[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(28[21:36])
    defparam i17577_2_lut.init = 16'h6666;
    LUT4 i17584_3_lut (.A(cnt_1mhz[2]), .B(cnt_1mhz[1]), .C(cnt_1mhz[0]), 
         .Z(n17[2])) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(28[21:36])
    defparam i17584_3_lut.init = 16'h6a6a;
    LUT4 i1_2_lut_3_lut_adj_27 (.A(\state_back_2__N_261[2] ), .B(n329), 
         .C(n331[17]), .Z(cnt_delay_19__N_187[17])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_27.init = 16'h2020;
    LUT4 i21355_2_lut_3_lut_4_lut (.A(cnt[1]), .B(n23114), .C(cnt[2]), 
         .D(cnt[0]), .Z(clk_c_enable_689)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i21355_2_lut_3_lut_4_lut.init = 16'h0020;
    LUT4 i17575_1_lut (.A(cnt_1mhz[0]), .Z(n17[0])) /* synthesis lut_function=(!(A)) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(28[21:36])
    defparam i17575_1_lut.init = 16'h5555;
    LUT4 data_wr_buffer_6__bdd_4_lut (.A(data_wr_buffer[6]), .B(cnt[2]), 
         .C(cnt[0]), .D(data_wr_buffer[7]), .Z(n24678)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;
    defparam data_wr_buffer_6__bdd_4_lut.init = 16'hfb0b;
    LUT4 i1376_1_lut (.A(cnt_init[0]), .Z(n1)) /* synthesis lut_function=(!(A)) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(100[21] 109[28])
    defparam i1376_1_lut.init = 16'h5555;
    LUT4 i3031_1_lut (.A(cnt_main[0]), .Z(n2_adj_5026)) /* synthesis lut_function=(!(A)) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(77[21] 95[28])
    defparam i3031_1_lut.init = 16'h5555;
    LUT4 i2629_3_lut (.A(\cnt_read[2] ), .B(cnt_read[1]), .C(cnt_read[0]), 
         .Z(n253[2])) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(142[48:63])
    defparam i2629_3_lut.init = 16'h6a6a;
    LUT4 i2622_2_lut (.A(cnt_read[1]), .B(cnt_read[0]), .Z(n253[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(142[48:63])
    defparam i2622_2_lut.init = 16'h6666;
    LUT4 i1_2_lut_adj_28 (.A(cnt_main[1]), .B(n23255), .Z(clk_c_enable_1422)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_28.init = 16'h8888;
    LUT4 n25707_bdd_4_lut (.A(n25707), .B(\state_back_2__N_261[2] ), .C(n25855), 
         .D(\state[1] ), .Z(n26776)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;
    defparam n25707_bdd_4_lut.init = 16'h11f0;
    LUT4 i21101_3_lut_4_lut_4_lut (.A(\state[1] ), .B(n25707), .C(\state[0] ), 
         .D(n25757), .Z(n23481)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(C (D)))) */ ;
    defparam i21101_3_lut_4_lut_4_lut.init = 16'h5808;
    LUT4 n329_bdd_3_lut_22217 (.A(n329), .B(n25757), .C(\state_back_2__N_261[2] ), 
         .Z(n25852)) /* synthesis lut_function=(A ((C)+!B)+!A !(B+(C))) */ ;
    defparam n329_bdd_3_lut_22217.init = 16'ha3a3;
    LUT4 n8345_bdd_4_lut (.A(n25669), .B(n25625), .C(n25741), .D(\state[0] ), 
         .Z(n25013)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B (C)+!B !((D)+!C)))) */ ;
    defparam n8345_bdd_4_lut.init = 16'h3faf;
    LUT4 i1_2_lut_3_lut_3_lut_4_lut_else_4_lut (.A(\state_back_2__N_261[2] ), 
         .B(n25680), .C(n25627), .D(n25592), .Z(n25775)) /* synthesis lut_function=(!(A (B+!(C))+!A (B+!(C (D))))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(44[14:19])
    defparam i1_2_lut_3_lut_3_lut_4_lut_else_4_lut.init = 16'h3020;
    LUT4 i13747_3_lut (.A(n5035), .B(cnt_write[1]), .C(cnt_write[0]), 
         .Z(cnt_write_3__N_333[1])) /* synthesis lut_function=(!(A+(B (C)+!B !(C)))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(115[30] 118[24])
    defparam i13747_3_lut.init = 16'h1414;
    LUT4 i1_2_lut_3_lut_adj_29 (.A(\state_back_2__N_261[2] ), .B(n329), 
         .C(n331[18]), .Z(cnt_delay_19__N_187[18])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_29.init = 16'h2020;
    CCU2D add_76_5 (.A0(cnt_delay[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt_delay[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n20480), .COUT(n20481), .S0(n331[3]), .S1(n331[4]));   // g:/fpga/mxo2/system/project/ds18b20z.v(161[43:59])
    defparam add_76_5.INIT0 = 16'h5aaa;
    defparam add_76_5.INIT1 = 16'h5aaa;
    defparam add_76_5.INJECT1_0 = "NO";
    defparam add_76_5.INJECT1_1 = "NO";
    CCU2D add_76_3 (.A0(cnt_delay[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt_delay[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n20479), .COUT(n20480), .S0(n331[1]), .S1(n331[2]));   // g:/fpga/mxo2/system/project/ds18b20z.v(161[43:59])
    defparam add_76_3.INIT0 = 16'h5aaa;
    defparam add_76_3.INIT1 = 16'h5aaa;
    defparam add_76_3.INJECT1_0 = "NO";
    defparam add_76_3.INJECT1_1 = "NO";
    PFUMX i22151 (.BLUT(n25766), .ALUT(n25767), .C0(\state_back_2__N_261[2] ), 
          .Z(num_delay_19__N_369[1]));
    LUT4 data_out_6__bdd_4_lut (.A(data_out[6]), .B(data_out[7]), .C(data_out[5]), 
         .D(tamp_out_11__N_414[1]), .Z(n1854[3])) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (B (C+(D))+!B !(C (D))))) */ ;
    defparam data_out_6__bdd_4_lut.init = 16'h1804;
    LUT4 data_wr_buffer_6__bdd_3_lut (.A(data_wr_buffer[4]), .B(cnt[2]), 
         .C(cnt[0]), .Z(n24679)) /* synthesis lut_function=(A (B+(C))) */ ;
    defparam data_wr_buffer_6__bdd_3_lut.init = 16'ha8a8;
    LUT4 i3392_3_lut_4_lut (.A(cnt[2]), .B(n25699), .C(n25705), .D(cnt_write[3]), 
         .Z(n5035)) /* synthesis lut_function=(A (B (D)+!B (C+(D)))+!A (C+(D))) */ ;
    defparam i3392_3_lut_4_lut.init = 16'hff70;
    LUT4 i21359_2_lut_3_lut_4_lut (.A(cnt[1]), .B(n23114), .C(cnt[2]), 
         .D(cnt[0]), .Z(clk_c_enable_557)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i21359_2_lut_3_lut_4_lut.init = 16'h0010;
    CCU2D sub_1360_add_2_21 (.A0(cnt_delay[19]), .B0(num_delay[12]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n20584), .S1(n329));
    defparam sub_1360_add_2_21.INIT0 = 16'h5999;
    defparam sub_1360_add_2_21.INIT1 = 16'h0000;
    defparam sub_1360_add_2_21.INJECT1_0 = "NO";
    defparam sub_1360_add_2_21.INJECT1_1 = "NO";
    LUT4 i21325_2_lut_3_lut_4_lut (.A(cnt[1]), .B(n23114), .C(cnt[2]), 
         .D(cnt[0]), .Z(clk_c_enable_1447)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i21325_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i28_3_lut (.A(cnt_init[0]), .B(\cnt_init[2] ), .C(cnt_init[1]), 
         .Z(n102[2])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(37[13:21])
    defparam i28_3_lut.init = 16'h6c6c;
    CCU2D sub_1360_add_2_19 (.A0(cnt_delay[17]), .B0(num_delay[12]), .C0(GND_net), 
          .D0(GND_net), .A1(cnt_delay[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n20583), .COUT(n20584));
    defparam sub_1360_add_2_19.INIT0 = 16'h5999;
    defparam sub_1360_add_2_19.INIT1 = 16'h5555;
    defparam sub_1360_add_2_19.INJECT1_0 = "NO";
    defparam sub_1360_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_1360_add_2_17 (.A0(cnt_delay[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt_delay[16]), .B1(num_delay[12]), .C1(GND_net), 
          .D1(GND_net), .CIN(n20582), .COUT(n20583));
    defparam sub_1360_add_2_17.INIT0 = 16'h5555;
    defparam sub_1360_add_2_17.INIT1 = 16'h5999;
    defparam sub_1360_add_2_17.INJECT1_0 = "NO";
    defparam sub_1360_add_2_17.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_adj_30 (.A(\state_back_2__N_261[2] ), .B(n329), 
         .C(n331[19]), .Z(cnt_delay_19__N_187[19])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_30.init = 16'h2020;
    LUT4 i21157_3_lut_4_lut (.A(cnt_init[1]), .B(n25707), .C(\state[0] ), 
         .D(n1853[0]), .Z(n2)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C)) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(100[21] 109[28])
    defparam i21157_3_lut_4_lut.init = 16'hf707;
    FD1P3AX state_i0_i2 (.D(state_2__N_258[2]), .SP(clk_c_enable_1371), 
            .CK(clk_c), .Q(\state_back_2__N_261[2] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam state_i0_i2.GSR = "ENABLED";
    FD1P3AX state_i0_i1 (.D(state_2__N_258[1]), .SP(clk_c_enable_1372), 
            .CK(clk_c), .Q(\state[1] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam state_i0_i1.GSR = "ENABLED";
    FD1P3AX cnt_read_i0_i0 (.D(n15869), .SP(clk_c_enable_1420), .CK(clk_c), 
            .Q(cnt_read[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam cnt_read_i0_i0.GSR = "ENABLED";
    FD1P3IX cnt_write_i0_i0 (.D(cnt_write_3__N_333[0]), .SP(clk_c_enable_1426), 
            .CD(n15328), .CK(clk_c), .Q(cnt_write[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam cnt_write_i0_i0.GSR = "ENABLED";
    LUT4 i12554_4_lut_then_2_lut (.A(\cnt_read[2] ), .B(cnt_read[1]), .Z(n25767)) /* synthesis lut_function=(!(A+(B))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(45[14:24])
    defparam i12554_4_lut_then_2_lut.init = 16'h1111;
    FD1S3IX cnt_1mhz_1980__i1 (.D(n17[1]), .CK(clk_c), .CD(n25765), .Q(cnt_1mhz[1]));   // g:/fpga/mxo2/system/project/ds18b20z.v(28[21:36])
    defparam cnt_1mhz_1980__i1.GSR = "ENABLED";
    FD1S3IX cnt_1mhz_1980__i2 (.D(n17[2]), .CK(clk_c), .CD(n25765), .Q(cnt_1mhz[2]));   // g:/fpga/mxo2/system/project/ds18b20z.v(28[21:36])
    defparam cnt_1mhz_1980__i2.GSR = "ENABLED";
    CCU2D sub_1360_add_2_15 (.A0(cnt_delay[13]), .B0(num_delay[12]), .C0(GND_net), 
          .D0(GND_net), .A1(cnt_delay[14]), .B1(num_delay[12]), .C1(GND_net), 
          .D1(GND_net), .CIN(n20581), .COUT(n20582));
    defparam sub_1360_add_2_15.INIT0 = 16'h5999;
    defparam sub_1360_add_2_15.INIT1 = 16'h5999;
    defparam sub_1360_add_2_15.INJECT1_0 = "NO";
    defparam sub_1360_add_2_15.INJECT1_1 = "NO";
    CCU2D add_76_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt_delay[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n20479), .S1(n331[0]));   // g:/fpga/mxo2/system/project/ds18b20z.v(161[43:59])
    defparam add_76_1.INIT0 = 16'hF000;
    defparam add_76_1.INIT1 = 16'h5555;
    defparam add_76_1.INJECT1_0 = "NO";
    defparam add_76_1.INJECT1_1 = "NO";
    CCU2D sub_1360_add_2_13 (.A0(cnt_delay[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt_delay[12]), .B1(num_delay[12]), .C1(GND_net), 
          .D1(GND_net), .CIN(n20580), .COUT(n20581));
    defparam sub_1360_add_2_13.INIT0 = 16'h5555;
    defparam sub_1360_add_2_13.INIT1 = 16'h5999;
    defparam sub_1360_add_2_13.INJECT1_0 = "NO";
    defparam sub_1360_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_1360_add_2_11 (.A0(cnt_delay[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt_delay[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n20579), .COUT(n20580));
    defparam sub_1360_add_2_11.INIT0 = 16'h5555;
    defparam sub_1360_add_2_11.INIT1 = 16'h5555;
    defparam sub_1360_add_2_11.INJECT1_0 = "NO";
    defparam sub_1360_add_2_11.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_31 (.A(cnt_main[3]), .B(cnt_main[0]), .C(cnt_main[2]), 
         .D(cnt_main[1]), .Z(n9)) /* synthesis lut_function=(!(A+(B (C (D))+!B !(D)))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam i1_4_lut_adj_31.init = 16'h1544;
    LUT4 i1_2_lut_adj_32 (.A(cnt_read[0]), .B(\cnt_read[2] ), .Z(n4)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_32.init = 16'h8888;
    CCU2D sub_1360_add_2_9 (.A0(cnt_delay[7]), .B0(num_delay[8]), .C0(GND_net), 
          .D0(GND_net), .A1(cnt_delay[8]), .B1(num_delay[8]), .C1(GND_net), 
          .D1(GND_net), .CIN(n20578), .COUT(n20579));
    defparam sub_1360_add_2_9.INIT0 = 16'h5999;
    defparam sub_1360_add_2_9.INIT1 = 16'h5999;
    defparam sub_1360_add_2_9.INJECT1_0 = "NO";
    defparam sub_1360_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_1360_add_2_7 (.A0(cnt_delay[5]), .B0(num_delay[5]), .C0(GND_net), 
          .D0(GND_net), .A1(cnt_delay[6]), .B1(num_delay[6]), .C1(GND_net), 
          .D1(GND_net), .CIN(n20577), .COUT(n20578));
    defparam sub_1360_add_2_7.INIT0 = 16'h5999;
    defparam sub_1360_add_2_7.INIT1 = 16'h5999;
    defparam sub_1360_add_2_7.INJECT1_0 = "NO";
    defparam sub_1360_add_2_7.INJECT1_1 = "NO";
    LUT4 i12554_4_lut_else_2_lut (.A(cnt_write[0]), .B(n25722), .C(cnt_write[1]), 
         .D(cnt_write[2]), .Z(n25766)) /* synthesis lut_function=(!(A ((D)+!B)+!A !(B (C+!(D))))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(45[14:24])
    defparam i12554_4_lut_else_2_lut.init = 16'h40cc;
    CCU2D sub_1360_add_2_5 (.A0(cnt_delay[3]), .B0(num_delay[3]), .C0(GND_net), 
          .D0(GND_net), .A1(cnt_delay[4]), .B1(num_delay[4]), .C1(GND_net), 
          .D1(GND_net), .CIN(n20576), .COUT(n20577));
    defparam sub_1360_add_2_5.INIT0 = 16'h5999;
    defparam sub_1360_add_2_5.INIT1 = 16'h5999;
    defparam sub_1360_add_2_5.INJECT1_0 = "NO";
    defparam sub_1360_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_1360_add_2_3 (.A0(cnt_delay[1]), .B0(num_delay[1]), .C0(GND_net), 
          .D0(GND_net), .A1(cnt_delay[2]), .B1(num_delay[2]), .C1(GND_net), 
          .D1(GND_net), .CIN(n20575), .COUT(n20576));
    defparam sub_1360_add_2_3.INIT0 = 16'h5999;
    defparam sub_1360_add_2_3.INIT1 = 16'h5999;
    defparam sub_1360_add_2_3.INJECT1_0 = "NO";
    defparam sub_1360_add_2_3.INJECT1_1 = "NO";
    LUT4 i13557_3_lut (.A(cnt[1]), .B(n20_adj_5027), .C(cnt[0]), .Z(cnt_2__N_161[1])) /* synthesis lut_function=(!(A (B+(C))+!A (B+!(C)))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(62[9] 163[16])
    defparam i13557_3_lut.init = 16'h1212;
    PFUMX i21642 (.BLUT(n24679), .ALUT(n24678), .C0(cnt[1]), .Z(one_wire_N_508));
    LUT4 i11848_3_lut_rep_302_4_lut (.A(cnt_write[3]), .B(n25668), .C(\state[0] ), 
         .D(n25669), .Z(n25584)) /* synthesis lut_function=(!(A (C+!(D))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(40[13:22])
    defparam i11848_3_lut_rep_302_4_lut.init = 16'h1f10;
    LUT4 one_wire_I_0_3_lut (.A(one_wire_out), .B(one_wire_N_505), .C(one_wire_N_510), 
         .Z(one_wire_N_504)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam one_wire_I_0_3_lut.init = 16'hcaca;
    LUT4 i3_4_lut (.A(one_wire_N_508), .B(cnt_write[2]), .C(n25663), .D(n25723), 
         .Z(one_wire_N_505)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i3_4_lut.init = 16'h2000;
    LUT4 i1_2_lut_rep_309_4_lut (.A(n25708), .B(\state_back_2__N_261[2] ), 
         .C(n25670), .D(n25680), .Z(n25591)) /* synthesis lut_function=(!(A (B+(D))+!A (B ((D)+!C)+!B (D)))) */ ;
    defparam i1_2_lut_rep_309_4_lut.init = 16'h0073;
    LUT4 i21504_2_lut_rep_405 (.A(\state_back_2__N_261[2] ), .B(\state[1] ), 
         .Z(n25687)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i21504_2_lut_rep_405.init = 16'h1111;
    LUT4 i1_2_lut_3_lut_adj_33 (.A(\state_back_2__N_261[2] ), .B(\state[1] ), 
         .C(n25757), .Z(n23372)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_33.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_34 (.A(\state_back_2__N_261[2] ), .B(\state[1] ), 
         .C(\state[0] ), .Z(n23154)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_34.init = 16'h1010;
    LUT4 i1_2_lut_rep_406 (.A(cnt_main[0]), .B(cnt_main[2]), .Z(n25688)) /* synthesis lut_function=(!((B)+!A)) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam i1_2_lut_rep_406.init = 16'h2222;
    LUT4 i1_2_lut_rep_344_3_lut_4_lut (.A(cnt_main[0]), .B(cnt_main[2]), 
         .C(cnt_main[3]), .D(cnt_main[1]), .Z(n25626)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam i1_2_lut_rep_344_3_lut_4_lut.init = 16'h0200;
    LUT4 i1_2_lut_rep_362_3_lut (.A(cnt_main[0]), .B(cnt_main[2]), .C(cnt_main[1]), 
         .Z(n25644)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam i1_2_lut_rep_362_3_lut.init = 16'h2020;
    LUT4 i13465_3_lut (.A(tamp_out_11__N_414[1]), .B(data_out[6]), .C(data_out[7]), 
         .Z(n1854[5])) /* synthesis lut_function=(A (B+(C))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(181[9] 201[16])
    defparam i13465_3_lut.init = 16'ha8a8;
    LUT4 i13016_3_lut_rep_407 (.A(\state[1] ), .B(\cnt_read[2] ), .C(\state_back_2__N_261[2] ), 
         .Z(n25689)) /* synthesis lut_function=(A (B (C))+!A (B+!(C))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(45[14:24])
    defparam i13016_3_lut_rep_407.init = 16'hc5c5;
    LUT4 i1_3_lut_4_lut_adj_35 (.A(\state[1] ), .B(\cnt_read[2] ), .C(\state_back_2__N_261[2] ), 
         .D(n3_adj_5028), .Z(num_delay_19__N_369[4])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(45[14:24])
    defparam i1_3_lut_4_lut_adj_35.init = 16'hcfc5;
    LUT4 i1_2_lut_3_lut_adj_36 (.A(cnt_write[0]), .B(cnt_write[1]), .C(cnt_write[2]), 
         .Z(n2_adj_5029)) /* synthesis lut_function=(A (C)+!A !(B+!(C))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(120[21] 134[28])
    defparam i1_2_lut_3_lut_adj_36.init = 16'hb0b0;
    LUT4 i3_4_lut_adj_37 (.A(n8250), .B(n23154), .C(cnt_main[3]), .D(n25618), 
         .Z(clk_c_enable_83)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam i3_4_lut_adj_37.init = 16'h0800;
    LUT4 i1_2_lut_adj_38 (.A(cnt_main[1]), .B(cnt_main[2]), .Z(n7_adj_5022)) /* synthesis lut_function=((B)+!A) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam i1_2_lut_adj_38.init = 16'hdddd;
    LUT4 i8_2_lut (.A(cnt_main[0]), .B(cnt_main[1]), .Z(n8250)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(34[13:21])
    defparam i8_2_lut.init = 16'h6666;
    LUT4 i21337_4_lut (.A(cnt_write[0]), .B(cnt_write[2]), .C(\state_back_2__N_261[2] ), 
         .D(n25618), .Z(n24052)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam i21337_4_lut.init = 16'h0100;
    LUT4 cnt_write_3__bdd_4_lut_22210 (.A(cnt_write[3]), .B(cnt_write[2]), 
         .C(cnt_write[0]), .D(cnt_write[1]), .Z(n25850)) /* synthesis lut_function=(A+(B ((D)+!C)+!B !(C+!(D)))) */ ;
    defparam cnt_write_3__bdd_4_lut_22210.init = 16'hefae;
    LUT4 tamp_out_11__N_414_1__bdd_4_lut_21660 (.A(tamp_out_11__N_414[1]), 
         .B(data_out[7]), .C(data_out[5]), .D(data_out[6]), .Z(n1854[2])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A !(B (C (D))+!B (D)))) */ ;
    defparam tamp_out_11__N_414_1__bdd_4_lut_21660.init = 16'h518a;
    LUT4 i1_2_lut_3_lut_adj_39 (.A(\state_back_2__N_261[2] ), .B(n329), 
         .C(n331[2]), .Z(cnt_delay_19__N_187[2])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_39.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_40 (.A(\state_back_2__N_261[2] ), .B(n329), 
         .C(n331[3]), .Z(cnt_delay_19__N_187[3])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_40.init = 16'h2020;
    LUT4 i21357_2_lut_2_lut_3_lut_4_lut (.A(cnt[0]), .B(cnt[2]), .C(n23114), 
         .D(cnt[1]), .Z(clk_c_enable_634)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i21357_2_lut_2_lut_3_lut_4_lut.init = 16'h0008;
    LUT4 i21353_2_lut_2_lut_3_lut_4_lut (.A(cnt[0]), .B(cnt[2]), .C(n23114), 
         .D(cnt[1]), .Z(clk_c_enable_747)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i21353_2_lut_2_lut_3_lut_4_lut.init = 16'h0800;
    LUT4 i13243_2_lut (.A(\cnt_read[2] ), .B(cnt_read[0]), .Z(n16018)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i13243_2_lut.init = 16'heeee;
    LUT4 tamp_out_11__N_414_1__bdd_4_lut_21936 (.A(tamp_out_11__N_414[1]), 
         .B(data_out[7]), .C(data_out[6]), .D(data_out[5]), .Z(n1854[1])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C (D)+!C !(D)))+!A (B ((D)+!C)+!B !(D)))) */ ;
    defparam tamp_out_11__N_414_1__bdd_4_lut_21936.init = 16'h3942;
    LUT4 i2_3_lut_adj_41 (.A(\state_back_2__N_261[2] ), .B(cnt_read[1]), 
         .C(\cnt_read[2] ), .Z(num_delay_19__N_369[0])) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i2_3_lut_adj_41.init = 16'h0808;
    LUT4 i21608_2_lut (.A(\state_back_2__N_261[2] ), .B(\state[1] ), .Z(n23827)) /* synthesis lut_function=(A+!(B)) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(62[9] 163[16])
    defparam i21608_2_lut.init = 16'hbbbb;
    LUT4 i2602_2_lut_rep_417 (.A(cnt[1]), .B(cnt[0]), .Z(n25699)) /* synthesis lut_function=(A (B)) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(138[77:87])
    defparam i2602_2_lut_rep_417.init = 16'h8888;
    LUT4 i2_2_lut_rep_370_3_lut (.A(cnt[1]), .B(cnt[0]), .C(cnt[2]), .Z(n25652)) /* synthesis lut_function=(A (B (C))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(138[77:87])
    defparam i2_2_lut_rep_370_3_lut.init = 16'h8080;
    LUT4 i13556_3_lut_4_lut (.A(cnt[1]), .B(cnt[0]), .C(n20_adj_5027), 
         .D(cnt[2]), .Z(cnt_2__N_161[2])) /* synthesis lut_function=(!(A (B (C+(D))+!B (C+!(D)))+!A (C+!(D)))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(138[77:87])
    defparam i13556_3_lut_4_lut.init = 16'h0708;
    FD1P3IX cnt_init_i0_i0 (.D(n1), .SP(clk_c_enable_1433), .CD(n12075), 
            .CK(clk_c), .Q(cnt_init[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam cnt_init_i0_i0.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_4_lut (.A(cnt[1]), .B(cnt[0]), .C(n25450), .D(cnt[2]), 
         .Z(n20_adj_5027)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(138[77:87])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hf8f0;
    LUT4 i2563_3_lut_4_lut (.A(cnt_main[1]), .B(cnt_main[0]), .C(cnt_main[2]), 
         .D(cnt_main[3]), .Z(n25[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;
    defparam i2563_3_lut_4_lut.init = 16'h7f80;
    LUT4 i2346_2_lut_3_lut (.A(cnt_main[1]), .B(cnt_main[0]), .C(cnt_main[2]), 
         .Z(n6)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i2346_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i2556_2_lut_3_lut (.A(cnt_main[1]), .B(cnt_main[0]), .C(cnt_main[2]), 
         .Z(n25[2])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;
    defparam i2556_2_lut_3_lut.init = 16'h7878;
    LUT4 tamp_out_11__N_414_1__bdd_4_lut (.A(tamp_out_11__N_414[1]), .B(data_out[7]), 
         .C(data_out[6]), .D(data_out[5]), .Z(n1854[4])) /* synthesis lut_function=(A (B (C (D))+!B !(C))+!A (B (C+(D)))) */ ;
    defparam tamp_out_11__N_414_1__bdd_4_lut.init = 16'hc642;
    FD1P3IX cnt_main_i0_i0 (.D(n2_adj_5026), .SP(clk_c_enable_1437), .CD(n14905), 
            .CK(clk_c), .Q(cnt_main[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam cnt_main_i0_i0.GSR = "ENABLED";
    FD1P3AX state_back_i0_i1 (.D(n25741), .SP(clk_c_enable_1416), .CK(clk_c), 
            .Q(state_back[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam state_back_i0_i1.GSR = "ENABLED";
    LUT4 i13931_3_lut_4_lut (.A(cnt_write[1]), .B(cnt_write[2]), .C(cnt_write[3]), 
         .D(cnt_write[0]), .Z(state_2__N_303[0])) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C (D))))) */ ;
    defparam i13931_3_lut_4_lut.init = 16'h0f1f;
    LUT4 i5_2_lut_rep_418 (.A(cnt_init[1]), .B(cnt_init[0]), .Z(n25700)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(37[13:21])
    defparam i5_2_lut_rep_418.init = 16'h6666;
    LUT4 i1_2_lut_3_lut_3_lut (.A(\cnt_init[2] ), .B(cnt_init[0]), .C(cnt_init[1]), 
         .Z(state_2__N_306[0])) /* synthesis lut_function=(!(A (B (C)+!B !(C)))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam i1_2_lut_3_lut_3_lut.init = 16'h7d7d;
    FD1P3IX cnt_read_i0_i2 (.D(n253[2]), .SP(clk_c_enable_1420), .CD(n12080), 
            .CK(clk_c), .Q(\cnt_read[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam cnt_read_i0_i2.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_adj_42 (.A(\state_back_2__N_261[2] ), .B(n329), 
         .C(n331[7]), .Z(cnt_delay_19__N_187[7])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_42.init = 16'h2020;
    FD1P3IX cnt_read_i0_i1 (.D(n253[1]), .SP(clk_c_enable_1420), .CD(n12080), 
            .CK(clk_c), .Q(cnt_read[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam cnt_read_i0_i1.GSR = "ENABLED";
    LUT4 i1_4_lut_4_lut (.A(\cnt_init[2] ), .B(\state[0] ), .C(n2_adj_5029), 
         .D(n25741), .Z(num_delay_19__N_369[6])) /* synthesis lut_function=(A (B (C (D)))+!A (B (C (D))+!B (D))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam i1_4_lut_4_lut.init = 16'hd100;
    LUT4 i21362_2_lut_3_lut_3_lut_4_lut (.A(cnt[2]), .B(cnt[0]), .C(cnt[1]), 
         .D(n23114), .Z(clk_c_enable_553)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i21362_2_lut_3_lut_3_lut_4_lut.init = 16'h0040;
    LUT4 i21368_2_lut_3_lut_3_lut_4_lut (.A(cnt[2]), .B(cnt[0]), .C(cnt[1]), 
         .D(n23114), .Z(clk_c_enable_201)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i21368_2_lut_3_lut_3_lut_4_lut.init = 16'h0004;
    LUT4 n25707_bdd_4_lut_22213 (.A(cnt_read[1]), .B(\state_back_2__N_261[2] ), 
         .C(\cnt_read[2] ), .D(cnt_read[0]), .Z(n25855)) /* synthesis lut_function=(A ((C+(D))+!B)+!A ((D)+!B)) */ ;
    defparam n25707_bdd_4_lut_22213.init = 16'hffb3;
    LUT4 i21541_4_lut_4_lut (.A(n25680), .B(n44), .C(n49), .D(n33), 
         .Z(clk_c_enable_1371)) /* synthesis lut_function=(!(A+(B (C+(D))+!B (C)))) */ ;
    defparam i21541_4_lut_4_lut.init = 16'h0105;
    LUT4 i4_4_lut (.A(n23656), .B(n23436), .C(\state_back_2__N_261[2] ), 
         .D(cnt_read[1]), .Z(n23114)) /* synthesis lut_function=((B+((D)+!C))+!A) */ ;
    defparam i4_4_lut.init = 16'hffdf;
    FD1P3AX temperature_i0_i8 (.D(temperature_buffer[0]), .SP(clk_c_enable_1422), 
            .CK(clk_c), .Q(temperature[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam temperature_i0_i8.GSR = "ENABLED";
    LUT4 i23_3_lut_4_lut_4_lut (.A(\state[0] ), .B(n25584), .C(\state[1] ), 
         .D(n25626), .Z(n32)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(62[9] 163[16])
    defparam i23_3_lut_4_lut_4_lut.init = 16'hcfc5;
    LUT4 i1_3_lut_3_lut (.A(\state[0] ), .B(\state[1] ), .C(n329), .Z(n33)) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(62[9] 163[16])
    defparam i1_3_lut_3_lut.init = 16'hcece;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut (.A(\state[0] ), .B(\state[1] ), .C(n25740), 
         .D(cnt_read[0]), .Z(n28)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(62[9] 163[16])
    defparam i1_2_lut_3_lut_4_lut_4_lut.init = 16'h0100;
    LUT4 state_2__I_0_216_Mux_0_i3_4_lut_4_lut (.A(\state[0] ), .B(n9), 
         .C(\state[1] ), .D(n2_adj_5024), .Z(n3_adj_5030)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A ((D)+!C)) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(62[9] 163[16])
    defparam state_2__I_0_216_Mux_0_i3_4_lut_4_lut.init = 16'hfd0d;
    LUT4 i3_4_lut_4_lut (.A(\state[0] ), .B(\cnt_init[2] ), .C(\state[1] ), 
         .D(cnt_init[0]), .Z(n21171)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(62[9] 163[16])
    defparam i3_4_lut_4_lut.init = 16'h1000;
    LUT4 i5600_2_lut_rep_310_3_lut_4_lut_4_lut (.A(\state[0] ), .B(cnt_main[3]), 
         .C(n25688), .D(cnt_main[1]), .Z(n25592)) /* synthesis lut_function=(!(A (B+!(C (D))))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(62[9] 163[16])
    defparam i5600_2_lut_rep_310_3_lut_4_lut_4_lut.init = 16'h7555;
    LUT4 i1_4_lut_4_lut_adj_43 (.A(\state[0] ), .B(cnt_main[3]), .C(clk_c_enable_1437), 
         .D(n6), .Z(n14905)) /* synthesis lut_function=(A (B (C (D)))+!A (C)) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(62[9] 163[16])
    defparam i1_4_lut_4_lut_adj_43.init = 16'hd050;
    LUT4 i18_4_lut_4_lut (.A(\state[0] ), .B(n23436), .C(\state_back_2__N_261[2] ), 
         .D(\cnt_read[2] ), .Z(n14)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C)+!B (C (D))))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(62[9] 163[16])
    defparam i18_4_lut_4_lut.init = 16'h0535;
    LUT4 i11_3_lut_4_lut_4_lut (.A(\state[0] ), .B(cnt_main[3]), .C(cnt_main[0]), 
         .D(cnt_main[1]), .Z(n14912)) /* synthesis lut_function=(!((B+(C (D)))+!A)) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(62[9] 163[16])
    defparam i11_3_lut_4_lut_4_lut.init = 16'h0222;
    LUT4 i1_4_lut_4_lut_adj_44 (.A(\state[0] ), .B(n15797), .C(\state[1] ), 
         .D(\state_back_2__N_261[2] ), .Z(num_delay_19__N_369[8])) /* synthesis lut_function=(!(A (C+(D))+!A (B (D)+!B (C+(D))))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(62[9] 163[16])
    defparam i1_4_lut_4_lut_adj_44.init = 16'h004f;
    LUT4 mux_83_Mux_2_i7_3_lut_4_lut (.A(cnt_read[1]), .B(\cnt_read[2] ), 
         .C(\state_back_2__N_261[2] ), .D(n21171), .Z(num_delay_19__N_369[2])) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(144[21] 155[28])
    defparam mux_83_Mux_2_i7_3_lut_4_lut.init = 16'hefe0;
    FD1P3IX cnt_write_i0_i3 (.D(cnt_write_3__N_333[3]), .SP(clk_c_enable_1426), 
            .CD(n15328), .CK(clk_c), .Q(cnt_write[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam cnt_write_i0_i3.GSR = "ENABLED";
    FD1P3IX cnt_write_i0_i2 (.D(cnt_write_3__N_333[2]), .SP(clk_c_enable_1426), 
            .CD(n15328), .CK(clk_c), .Q(cnt_write[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam cnt_write_i0_i2.GSR = "ENABLED";
    LUT4 i2364_2_lut_rep_423 (.A(cnt_write[1]), .B(cnt_write[2]), .Z(n25705)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2364_2_lut_rep_423.init = 16'h8888;
    LUT4 i1_3_lut_4_lut_3_lut (.A(cnt_write[1]), .B(cnt_write[2]), .C(cnt_write[0]), 
         .Z(n34)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;
    defparam i1_3_lut_4_lut_3_lut.init = 16'h8e8e;
    LUT4 i2345_2_lut_rep_373_3_lut (.A(cnt_write[1]), .B(cnt_write[2]), 
         .C(cnt_write[3]), .Z(n25655)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i2345_2_lut_rep_373_3_lut.init = 16'hf8f8;
    LUT4 i21341_2_lut_rep_425 (.A(cnt_init[0]), .B(\cnt_init[2] ), .Z(n25707)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i21341_2_lut_rep_425.init = 16'h1111;
    LUT4 i85_4_lut_3_lut (.A(cnt_init[0]), .B(\cnt_init[2] ), .C(cnt_init[1]), 
         .Z(n16451)) /* synthesis lut_function=((B (C))+!A) */ ;
    defparam i85_4_lut_3_lut.init = 16'hd5d5;
    LUT4 i1_2_lut_rep_397_3_lut (.A(cnt_init[0]), .B(\cnt_init[2] ), .C(\state[1] ), 
         .Z(n25679)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_rep_397_3_lut.init = 16'h1010;
    FD1P3IX cnt_write_i0_i1 (.D(cnt_write_3__N_333[1]), .SP(clk_c_enable_1426), 
            .CD(n15328), .CK(clk_c), .Q(cnt_write[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam cnt_write_i0_i1.GSR = "ENABLED";
    LUT4 i21499_2_lut (.A(cnt[0]), .B(n20_adj_5027), .Z(cnt_2__N_161[0])) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i21499_2_lut.init = 16'h1111;
    LUT4 i1_2_lut_rep_426 (.A(\state[0] ), .B(\state[1] ), .Z(n25708)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_426.init = 16'heeee;
    LUT4 i21470_2_lut_2_lut_3_lut_4_lut (.A(\state[0] ), .B(\state[1] ), 
         .C(n25765), .D(clk_1mhz), .Z(clk_c_enable_1420)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i21470_2_lut_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i1_2_lut_3_lut_adj_45 (.A(\state[0] ), .B(\state[1] ), .C(cnt_read[0]), 
         .Z(n23436)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_3_lut_adj_45.init = 16'hfefe;
    LUT4 n5035_bdd_3_lut_22089_4_lut (.A(\state[0] ), .B(\state[1] ), .C(\cnt_read[2] ), 
         .D(n23814), .Z(n25451)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam n5035_bdd_3_lut_22089_4_lut.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_adj_46 (.A(\state[0] ), .B(\state[1] ), .C(cnt_read[1]), 
         .Z(n4_adj_5025)) /* synthesis lut_function=(A+(B+!(C))) */ ;
    defparam i1_2_lut_3_lut_adj_46.init = 16'hefef;
    LUT4 i20762_2_lut (.A(cnt_init[1]), .B(\state[0] ), .Z(n23622)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i20762_2_lut.init = 16'heeee;
    CCU2D sub_1360_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt_delay[0]), .B1(num_delay[0]), .C1(GND_net), 
          .D1(GND_net), .COUT(n20575));
    defparam sub_1360_add_2_1.INIT0 = 16'h0000;
    defparam sub_1360_add_2_1.INIT1 = 16'h5999;
    defparam sub_1360_add_2_1.INJECT1_0 = "NO";
    defparam sub_1360_add_2_1.INJECT1_1 = "NO";
    LUT4 i21338_3_lut_4_lut (.A(cnt_write[1]), .B(cnt_write[3]), .C(n24052), 
         .D(n25722), .Z(clk_c_enable_86)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i21338_3_lut_4_lut.init = 16'h1000;
    LUT4 i2_3_lut_4_lut (.A(cnt_write[1]), .B(cnt_write[3]), .C(cnt_write[2]), 
         .D(cnt_write[0]), .Z(n1853[0])) /* synthesis lut_function=(A+(B+!(C (D)))) */ ;
    defparam i2_3_lut_4_lut.init = 16'hefff;
    LUT4 i1_2_lut_rep_435 (.A(cnt_main[1]), .B(cnt_main[2]), .Z(n25717)) /* synthesis lut_function=(A (B)) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam i1_2_lut_rep_435.init = 16'h8888;
    LUT4 i13920_1_lut_2_lut (.A(cnt_main[1]), .B(cnt_main[2]), .Z(n7_adj_5023)) /* synthesis lut_function=(!(A (B))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam i13920_1_lut_2_lut.init = 16'h7777;
    LUT4 i2_4_lut_4_lut (.A(n25741), .B(n46), .C(n25627), .D(n50), .Z(clk_c_enable_683)) /* synthesis lut_function=(A (B (C (D)))+!A (C (D))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(44[14:19])
    defparam i2_4_lut_4_lut.init = 16'hd000;
    LUT4 i1_2_lut_3_lut_3_lut_4_lut_then_4_lut (.A(\state_back_2__N_261[2] ), 
         .B(n25584), .C(n25680), .D(n25627), .Z(n25776)) /* synthesis lut_function=(!(A (C+!(D))+!A ((C+!(D))+!B))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(44[14:19])
    defparam i1_2_lut_3_lut_3_lut_4_lut_then_4_lut.init = 16'h0e00;
    LUT4 i1_2_lut_adj_47 (.A(\cnt_init[2] ), .B(cnt_init[1]), .Z(n15797)) /* synthesis lut_function=(A+!(B)) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam i1_2_lut_adj_47.init = 16'hbbbb;
    LUT4 i2806_3_lut_4_lut (.A(cnt_write[0]), .B(cnt_write[1]), .C(n5035), 
         .D(cnt_write[2]), .Z(cnt_write_3__N_333[3])) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(115[30] 118[24])
    defparam i2806_3_lut_4_lut.init = 16'h0800;
    LUT4 i1_2_lut_rep_441 (.A(cnt_write[0]), .B(cnt_write[1]), .Z(n25723)) /* synthesis lut_function=(A (B)) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(115[30] 118[24])
    defparam i1_2_lut_rep_441.init = 16'h8888;
    LUT4 i13817_2_lut_3_lut_4_lut (.A(\state[1] ), .B(\state[0] ), .C(n25668), 
         .D(cnt_write[3]), .Z(n16602)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i13817_2_lut_3_lut_4_lut.init = 16'h8880;
    LUT4 i4_4_lut_adj_48 (.A(\cnt_init[2] ), .B(cnt_init[0]), .C(one_wire_out), 
         .D(n23622), .Z(n21141)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i4_4_lut_adj_48.init = 16'h0002;
    LUT4 i20874_2_lut_rep_440 (.A(\state[1] ), .B(\state[0] ), .Z(n25722)) /* synthesis lut_function=(A (B)) */ ;
    defparam i20874_2_lut_rep_440.init = 16'h8888;
    LUT4 i2_3_lut_rep_381_4_lut (.A(\state[1] ), .B(\state[0] ), .C(\state_back_2__N_261[2] ), 
         .D(cnt_write[3]), .Z(n25663)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i2_3_lut_rep_381_4_lut.init = 16'h0008;
    LUT4 i1_2_lut_3_lut_adj_49 (.A(\state_back_2__N_261[2] ), .B(n329), 
         .C(n331[4]), .Z(cnt_delay_19__N_187[4])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_49.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_50 (.A(\state_back_2__N_261[2] ), .B(n329), 
         .C(n331[8]), .Z(cnt_delay_19__N_187[8])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_50.init = 16'h2020;
    LUT4 i5335_2_lut_rep_456 (.A(cnt_write[0]), .B(cnt_write[1]), .Z(n25738)) /* synthesis lut_function=(A+!(B)) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(120[21] 134[28])
    defparam i5335_2_lut_rep_456.init = 16'hbbbb;
    LUT4 i11819_3_lut_rep_386_4_lut_3_lut (.A(cnt_write[0]), .B(cnt_write[1]), 
         .C(cnt_write[2]), .Z(n25668)) /* synthesis lut_function=(!(A (B (C))+!A (B+(C)))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(120[21] 134[28])
    defparam i11819_3_lut_rep_386_4_lut_3_lut.init = 16'h2b2b;
    LUT4 i1_2_lut_rep_457 (.A(\cnt_init[2] ), .B(cnt_init[1]), .Z(n25739)) /* synthesis lut_function=(A (B)) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam i1_2_lut_rep_457.init = 16'h8888;
    LUT4 i1_2_lut_rep_387_3_lut (.A(\cnt_init[2] ), .B(cnt_init[1]), .C(cnt_init[0]), 
         .Z(n25669)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam i1_2_lut_rep_387_3_lut.init = 16'h7070;
    CCU2D add_76_21 (.A0(cnt_delay[19]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n20488), 
          .S0(n331[19]));   // g:/fpga/mxo2/system/project/ds18b20z.v(161[43:59])
    defparam add_76_21.INIT0 = 16'h5aaa;
    defparam add_76_21.INIT1 = 16'h0000;
    defparam add_76_21.INJECT1_0 = "NO";
    defparam add_76_21.INJECT1_1 = "NO";
    LUT4 i13375_2_lut_rep_458 (.A(cnt_read[1]), .B(\cnt_read[2] ), .Z(n25740)) /* synthesis lut_function=(A (B)) */ ;
    defparam i13375_2_lut_rep_458.init = 16'h8888;
    LUT4 i13563_2_lut_rep_388_3_lut (.A(cnt_read[1]), .B(\cnt_read[2] ), 
         .C(cnt_read[0]), .Z(n25670)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13563_2_lut_rep_388_3_lut.init = 16'h7070;
    LUT4 i1_2_lut_rep_331_3_lut_3_lut_4_lut (.A(cnt_read[1]), .B(\cnt_read[2] ), 
         .C(cnt_read[0]), .D(\state[0] ), .Z(n25613)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A ((D)+!C))) */ ;
    defparam i1_2_lut_rep_331_3_lut_3_lut_4_lut.init = 16'h0070;
    LUT4 i21546_2_lut_rep_459 (.A(\state[1] ), .B(\state_back_2__N_261[2] ), 
         .Z(n25741)) /* synthesis lut_function=(!((B)+!A)) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(44[14:19])
    defparam i21546_2_lut_rep_459.init = 16'h2222;
    LUT4 i8897_2_lut_rep_460 (.A(\state[0] ), .B(\state[1] ), .Z(n25742)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i8897_2_lut_rep_460.init = 16'hbbbb;
    LUT4 i1_2_lut_3_lut_adj_51 (.A(\state[0] ), .B(\state[1] ), .C(\state_back_2__N_261[2] ), 
         .Z(state_back_2__N_261[0])) /* synthesis lut_function=(!(A (C)+!A (B+(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_51.init = 16'h0b0b;
    CCU2D add_76_11 (.A0(cnt_delay[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt_delay[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n20483), .COUT(n20484), .S0(n331[9]), .S1(n331[10]));   // g:/fpga/mxo2/system/project/ds18b20z.v(161[43:59])
    defparam add_76_11.INIT0 = 16'h5aaa;
    defparam add_76_11.INIT1 = 16'h5aaa;
    defparam add_76_11.INJECT1_0 = "NO";
    defparam add_76_11.INJECT1_1 = "NO";
    LUT4 i2929_1_lut (.A(one_wire_N_502), .Z(n5709)) /* synthesis lut_function=(!(A)) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(48[1] 165[4])
    defparam i2929_1_lut.init = 16'h5555;
    FD1P3IX cnt_init_i0_i2 (.D(n102[2]), .SP(clk_c_enable_1433), .CD(n12075), 
            .CK(clk_c), .Q(\cnt_init[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam cnt_init_i0_i2.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_adj_52 (.A(\state_back_2__N_261[2] ), .B(n329), 
         .C(n331[0]), .Z(n23294)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_52.init = 16'h2020;
    LUT4 n14645_bdd_2_lut_4_lut (.A(n25669), .B(n25625), .C(\state[0] ), 
         .D(\state_back_2__N_261[2] ), .Z(n25482)) /* synthesis lut_function=(!(A (B (C+(D))+!B (D))+!A (B+((D)+!C)))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(44[14:19])
    defparam n14645_bdd_2_lut_4_lut.init = 16'h003a;
    LUT4 i1_2_lut_4_lut_adj_53 (.A(n25669), .B(n25625), .C(\state[0] ), 
         .D(\state[1] ), .Z(n37)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B (D)+!B !(C+!(D))))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(44[14:19])
    defparam i1_2_lut_4_lut_adj_53.init = 16'h3aff;
    LUT4 i1_2_lut_adj_54 (.A(cnt_main[1]), .B(n23255), .Z(clk_c_enable_709)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut_adj_54.init = 16'h4444;
    LUT4 i2_4_lut (.A(clk_c_enable_1437), .B(\state[0] ), .C(n66), .D(cnt_main[3]), 
         .Z(n23255)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i2_4_lut.init = 16'h0800;
    LUT4 i1_2_lut_adj_55 (.A(cnt_main[0]), .B(cnt_main[2]), .Z(n66)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_55.init = 16'heeee;
    LUT4 i49_4_lut (.A(n25669), .B(cnt_write[3]), .C(\state[0] ), .D(n34), 
         .Z(n46)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B+!(C (D))))) */ ;
    defparam i49_4_lut.init = 16'h3a0a;
    LUT4 n14645_bdd_3_lut_4_lut (.A(\state[0] ), .B(n25626), .C(\state_back_2__N_261[2] ), 
         .D(n25613), .Z(n25483)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam n14645_bdd_3_lut_4_lut.init = 16'hf808;
    FD1P3IX cnt_init_i0_i1 (.D(n25700), .SP(clk_c_enable_1433), .CD(n12075), 
            .CK(clk_c), .Q(cnt_init[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam cnt_init_i0_i1.GSR = "ENABLED";
    FD1P3IX cnt_main_i0_i3 (.D(n25[3]), .SP(clk_c_enable_1437), .CD(n14905), 
            .CK(clk_c), .Q(cnt_main[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam cnt_main_i0_i3.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_343_4_lut_4_lut (.A(cnt_write[0]), .B(cnt_write[1]), 
         .C(cnt_write[2]), .D(cnt_write[3]), .Z(n25625)) /* synthesis lut_function=(A (((D)+!C)+!B)+!A (B (D)+!B ((D)+!C))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(40[13:22])
    defparam i1_2_lut_rep_343_4_lut_4_lut.init = 16'hff2b;
    LUT4 i1_2_lut_3_lut_adj_56 (.A(\state_back_2__N_261[2] ), .B(n329), 
         .C(n331[10]), .Z(cnt_delay_19__N_187[10])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_56.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_57 (.A(\state_back_2__N_261[2] ), .B(n329), 
         .C(n331[1]), .Z(cnt_delay_19__N_187[1])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_57.init = 16'h2020;
    LUT4 i3_4_lut_adj_58 (.A(cnt_main[3]), .B(n23154), .C(n25680), .D(n25644), 
         .Z(clk_c_enable_717)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i3_4_lut_adj_58.init = 16'h0800;
    LUT4 i1_2_lut_adj_59 (.A(\state[1] ), .B(n46), .Z(n29)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i1_2_lut_adj_59.init = 16'hdddd;
    PFUMX i22104 (.BLUT(n25483), .ALUT(n25482), .C0(\state[1] ), .Z(n25484));
    LUT4 i13028_4_lut (.A(n15797), .B(cnt_write[2]), .C(\state[0] ), .D(n25738), 
         .Z(n3_adj_5028)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(44[14:19])
    defparam i13028_4_lut.init = 16'hca0a;
    LUT4 i9122_2_lut (.A(\cnt_read[2] ), .B(\state_back_2__N_261[2] ), .Z(num_delay_19__N_369[3])) /* synthesis lut_function=(A (B)) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(62[9] 163[16])
    defparam i9122_2_lut.init = 16'h8888;
    CCU2D add_76_9 (.A0(cnt_delay[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt_delay[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n20482), .COUT(n20483), .S0(n331[7]), .S1(n331[8]));   // g:/fpga/mxo2/system/project/ds18b20z.v(161[43:59])
    defparam add_76_9.INIT0 = 16'h5aaa;
    defparam add_76_9.INIT1 = 16'h5aaa;
    defparam add_76_9.INJECT1_0 = "NO";
    defparam add_76_9.INJECT1_1 = "NO";
    PFUMX i22102 (.BLUT(n25480), .ALUT(n25475), .C0(\state_back_2__N_261[2] ), 
          .Z(state_2__N_258[2]));
    PFUMX i22100 (.BLUT(n25477), .ALUT(n25476), .C0(\state[1] ), .Z(n25478));
    CCU2D add_76_19 (.A0(cnt_delay[17]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt_delay[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n20487), .COUT(n20488), .S0(n331[17]), .S1(n331[18]));   // g:/fpga/mxo2/system/project/ds18b20z.v(161[43:59])
    defparam add_76_19.INIT0 = 16'h5aaa;
    defparam add_76_19.INIT1 = 16'h5aaa;
    defparam add_76_19.INJECT1_0 = "NO";
    defparam add_76_19.INJECT1_1 = "NO";
    CCU2D add_76_13 (.A0(cnt_delay[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt_delay[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n20484), .COUT(n20485), .S0(n331[11]), .S1(n331[12]));   // g:/fpga/mxo2/system/project/ds18b20z.v(161[43:59])
    defparam add_76_13.INIT0 = 16'h5aaa;
    defparam add_76_13.INIT1 = 16'h5aaa;
    defparam add_76_13.INJECT1_0 = "NO";
    defparam add_76_13.INJECT1_1 = "NO";
    CCU2D add_76_17 (.A0(cnt_delay[15]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt_delay[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n20486), .COUT(n20487), .S0(n331[15]), .S1(n331[16]));   // g:/fpga/mxo2/system/project/ds18b20z.v(161[43:59])
    defparam add_76_17.INIT0 = 16'h5aaa;
    defparam add_76_17.INIT1 = 16'h5aaa;
    defparam add_76_17.INJECT1_0 = "NO";
    defparam add_76_17.INJECT1_1 = "NO";
    LUT4 i2_4_lut_adj_60 (.A(clk_1mhz), .B(n25765), .C(n24036), .D(\state[1] ), 
         .Z(clk_c_enable_736)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i2_4_lut_adj_60.init = 16'h0004;
    CCU2D add_76_15 (.A0(cnt_delay[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt_delay[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n20485), .COUT(n20486), .S0(n331[13]), .S1(n331[14]));   // g:/fpga/mxo2/system/project/ds18b20z.v(161[43:59])
    defparam add_76_15.INIT0 = 16'h5aaa;
    defparam add_76_15.INIT1 = 16'h5aaa;
    defparam add_76_15.INJECT1_0 = "NO";
    defparam add_76_15.INJECT1_1 = "NO";
    LUT4 i21321_2_lut (.A(\state_back_2__N_261[2] ), .B(\state[0] ), .Z(n24036)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i21321_2_lut.init = 16'h6666;
    LUT4 i2_3_lut_rep_475 (.A(cnt_main[0]), .B(cnt_main[3]), .C(cnt_main[2]), 
         .Z(n25757)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;
    defparam i2_3_lut_rep_475.init = 16'h0404;
    PFUMX i22090 (.BLUT(n25452), .ALUT(n25451), .C0(\state_back_2__N_261[2] ), 
          .Z(n25453));
    LUT4 i1_2_lut_3_lut_adj_61 (.A(\state_back_2__N_261[2] ), .B(n329), 
         .C(n331[5]), .Z(cnt_delay_19__N_187[5])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_61.init = 16'h2020;
    FD1P3IX cnt_main_i0_i2 (.D(n25[2]), .SP(clk_c_enable_1437), .CD(n14905), 
            .CK(clk_c), .Q(cnt_main[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam cnt_main_i0_i2.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_adj_62 (.A(\state_back_2__N_261[2] ), .B(n329), 
         .C(n331[11]), .Z(cnt_delay_19__N_187[11])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_62.init = 16'h2020;
    LUT4 i2348_3_lut_rep_483 (.A(cnt_1mhz[0]), .B(cnt_1mhz[2]), .C(cnt_1mhz[1]), 
         .Z(n25765)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i2348_3_lut_rep_483.init = 16'hc8c8;
    PFUMX i22087 (.BLUT(n25449), .ALUT(n25448), .C0(\state_back_2__N_261[2] ), 
          .Z(n25450));
    LUT4 i97_2_lut_rep_398_4_lut (.A(cnt_1mhz[0]), .B(cnt_1mhz[2]), .C(cnt_1mhz[1]), 
         .D(clk_1mhz), .Z(n25680)) /* synthesis lut_function=(A ((D)+!B)+!A (((D)+!C)+!B)) */ ;
    defparam i97_2_lut_rep_398_4_lut.init = 16'hff37;
    LUT4 clk_1mhz_I_0_2_lut_4_lut (.A(cnt_1mhz[0]), .B(cnt_1mhz[2]), .C(cnt_1mhz[1]), 
         .D(clk_1mhz), .Z(clk_1mhz_N_503)) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A (B (C (D)+!C !(D))+!B !(D)))) */ ;
    defparam clk_1mhz_I_0_2_lut_4_lut.init = 16'h37c8;
    LUT4 i1_2_lut_3_lut_adj_63 (.A(\state_back_2__N_261[2] ), .B(n329), 
         .C(n331[9]), .Z(cnt_delay_19__N_187[9])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_63.init = 16'h2020;
    PFUMX i12 (.BLUT(n3_adj_5030), .ALUT(n7), .C0(\state_back_2__N_261[2] ), 
          .Z(state_2__N_258[0]));
    FD1P3IX cnt_main_i0_i1 (.D(n8250), .SP(clk_c_enable_1437), .CD(n14905), 
            .CK(clk_c), .Q(cnt_main[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam cnt_main_i0_i1.GSR = "ENABLED";
    FD1P3AX cnt_i0_i2 (.D(cnt_2__N_161[2]), .SP(clk_c_enable_1439), .CK(clk_c), 
            .Q(cnt[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam cnt_i0_i2.GSR = "ENABLED";
    FD1P3AX cnt_i0_i1 (.D(cnt_2__N_161[1]), .SP(clk_c_enable_1439), .CK(clk_c), 
            .Q(cnt[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam cnt_i0_i1.GSR = "ENABLED";
    PFUMX i54 (.BLUT(n30), .ALUT(n23372), .C0(\state[0] ), .Z(n49));
    FD1P3AX temperature_buffer_i0_i0 (.D(one_wire_out), .SP(clk_c_enable_1447), 
            .CK(clk_c), .Q(temperature_buffer[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=61, LSE_RLINE=67 */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(61[14] 164[8])
    defparam temperature_buffer_i0_i0.GSR = "DISABLED";
    LUT4 i17_4_lut_adj_64 (.A(n25707), .B(cnt_write[0]), .C(\state[0] ), 
         .D(n25655), .Z(n13)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // g:/fpga/mxo2/system/project/ds18b20z.v(44[14:19])
    defparam i17_4_lut_adj_64.init = 16'h0aca;
    L6MUX21 i22208 (.D0(n26776), .D1(n25853), .SD(\state[0] ), .Z(n25857));
    LUT4 i20937_3_lut_4_lut (.A(cnt[2]), .B(n25699), .C(cnt_read[0]), 
         .D(cnt_read[1]), .Z(n23814)) /* synthesis lut_function=(A (B (D)+!B (C+(D)))+!A (C+(D))) */ ;
    defparam i20937_3_lut_4_lut.init = 16'hff70;
    
endmodule
